magic
tech sky130A
timestamp 1697774992
<< poly >>
rect 2590 7245 2620 7260
rect 1480 5860 1515 5875
rect 1480 5790 1495 5860
rect 1455 5775 1495 5790
rect 1445 4435 1500 4450
rect 1485 3180 1500 4435
rect 1485 3165 1525 3180
<< locali >>
rect 2590 7190 2620 7215
rect 1445 5710 1495 5730
rect 1475 4605 1495 5710
rect 1475 4560 1525 4605
rect 1470 4490 1530 4510
rect 1470 4420 1490 4490
rect 2595 4480 2620 4510
<< metal1 >>
rect -280 7105 -265 8295
rect -280 4500 -265 6995
rect 1500 5920 1515 7110
rect 2605 5920 2620 7110
rect 1500 4625 1515 5815
rect 2605 4625 2620 5815
rect -280 3205 -265 4385
rect 1500 3240 1515 4430
rect 2605 3240 2620 4430
use diff_amp  diff_amp_0
timestamp 1697719741
transform 1 0 2230 0 1 3220
box -730 -55 390 4040
use v_gen  v_gen_0
timestamp 1697774992
transform 1 0 -10 0 1 5660
box -270 -2540 1480 2675
<< labels >>
rlabel poly 2620 7250 2620 7250 3 Vref
rlabel metal1 1500 5220 1500 5220 7 VP
rlabel metal1 1500 6515 1500 6515 7 VN
rlabel locali 2620 7205 2620 7205 3 Vin
rlabel metal1 -280 3795 -280 3795 7 VP
rlabel locali 2620 4495 2620 4495 7 Vout
rlabel metal1 -280 7710 -280 7710 7 VP
rlabel locali 1500 4500 1500 4500 7 Vbp
rlabel metal1 -280 5744 -280 5744 7 VN
rlabel locali 1500 4570 1500 4570 7 Vcp
rlabel metal1 1500 3830 1500 3830 7 VN
<< end >>
