magic
tech sky130A
timestamp 1694522166
<< nwell >>
rect -120 130 150 270
<< nmos >>
rect 0 -5 15 95
rect 65 -5 80 95
<< pmos >>
rect 0 150 15 250
rect 65 150 80 250
<< ndiff >>
rect -50 80 0 95
rect -50 10 -35 80
rect -15 10 0 80
rect -50 -5 0 10
rect 15 80 65 95
rect 15 10 30 80
rect 50 10 65 80
rect 15 -5 65 10
rect 80 80 130 95
rect 80 10 95 80
rect 115 10 130 80
rect 80 -5 130 10
<< pdiff >>
rect -50 235 0 250
rect -50 165 -35 235
rect -15 165 0 235
rect -50 150 0 165
rect 15 235 65 250
rect 15 165 30 235
rect 50 165 65 235
rect 15 150 65 165
rect 80 235 130 250
rect 80 165 95 235
rect 115 165 130 235
rect 80 150 130 165
<< ndiffc >>
rect -35 10 -15 80
rect 30 10 50 80
rect 95 10 115 80
<< pdiffc >>
rect -35 165 -15 235
rect 30 165 50 235
rect 95 165 115 235
<< psubdiff >>
rect -100 80 -50 95
rect -100 10 -85 80
rect -65 10 -50 80
rect -100 -5 -50 10
<< nsubdiff >>
rect -100 235 -50 250
rect -100 165 -85 235
rect -65 165 -50 235
rect -100 150 -50 165
<< psubdiffcont >>
rect -85 10 -65 80
<< nsubdiffcont >>
rect -85 165 -65 235
<< poly >>
rect 0 250 15 265
rect 65 250 80 265
rect 0 95 15 150
rect 65 95 80 150
rect 0 -20 15 -5
rect 65 -20 80 -5
rect -25 -30 15 -20
rect -25 -50 -15 -30
rect 5 -50 15 -30
rect -25 -60 15 -50
rect 40 -30 80 -20
rect 40 -50 50 -30
rect 70 -50 80 -30
rect 40 -60 80 -50
<< polycont >>
rect -15 -50 5 -30
rect 50 -50 70 -30
<< locali >>
rect -95 235 -5 245
rect -95 165 -85 235
rect -65 165 -35 235
rect -15 165 -5 235
rect -95 155 -5 165
rect 20 235 60 245
rect 20 165 30 235
rect 50 165 60 235
rect 20 155 60 165
rect 85 235 125 245
rect 85 165 95 235
rect 115 165 125 235
rect 85 155 125 165
rect 40 130 60 155
rect 40 110 105 130
rect 85 90 105 110
rect -95 80 -5 90
rect -95 10 -85 80
rect -65 10 -35 80
rect -15 10 -5 80
rect -95 0 -5 10
rect 20 80 60 90
rect 20 10 30 80
rect 50 10 60 80
rect 20 0 60 10
rect 85 80 125 90
rect 85 10 95 80
rect 115 10 125 80
rect 85 0 125 10
rect 105 -20 125 0
rect -120 -30 15 -20
rect -120 -40 -15 -30
rect -25 -50 -15 -40
rect 5 -50 15 -30
rect -25 -60 15 -50
rect 40 -30 80 -20
rect 40 -50 50 -30
rect 70 -50 80 -30
rect 105 -40 150 -20
rect 40 -60 80 -50
rect 40 -80 60 -60
rect -120 -100 60 -80
<< viali >>
rect -85 165 -65 235
rect -35 165 -15 235
rect 95 165 115 235
rect -85 10 -65 80
rect -35 10 -15 80
<< metal1 >>
rect -120 235 150 245
rect -120 165 -85 235
rect -65 165 -35 235
rect -15 165 95 235
rect 115 165 150 235
rect -120 155 150 165
rect -120 80 150 90
rect -120 10 -85 80
rect -65 10 -35 80
rect -15 10 150 80
rect -120 0 150 10
<< labels >>
rlabel locali 150 -30 150 -30 3 Y
port 3 e
rlabel metal1 -120 45 -120 45 7 VN
port 5 w
rlabel metal1 -120 200 -120 200 7 VP
port 4 w
rlabel locali -120 -90 -120 -90 7 A
port 1 w
rlabel locali -120 -30 -120 -30 7 B
port 2 w
<< end >>
