* SPICE3 file created from buffer.ext - technology: sky130A

.subckt inverter A Y VN VP
X0 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

.subckt buffer
Xinverter_0 A inverter_1/A VN VP inverter
Xinverter_1 inverter_1/A Y VN VP inverter
.ends

