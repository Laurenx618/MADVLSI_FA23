magic
tech sky130A
timestamp 1698134288
<< nwell >>
rect -370 1420 1580 2670
rect -370 -2520 1580 -1280
<< nmos >>
rect -300 140 -250 1340
rect -200 140 -150 1340
rect 30 140 80 1340
rect 130 140 180 1340
rect 230 140 280 1340
rect 330 140 380 1340
rect 430 140 480 1340
rect 530 140 580 1340
rect 630 140 680 1340
rect 730 140 780 1340
rect 830 140 880 1340
rect 930 140 980 1340
rect 1030 140 1080 1340
rect 1130 140 1180 1340
rect 1360 140 1410 1340
rect 1460 140 1510 1340
rect -300 -1200 -250 0
rect -200 -1200 -150 0
rect 30 -1200 80 0
rect 130 -1200 180 0
rect 230 -1200 280 0
rect 330 -1200 380 0
rect 430 -1200 480 0
rect 530 -1200 580 0
rect 630 -1200 680 0
rect 730 -1200 780 0
rect 830 -1200 880 0
rect 930 -1200 980 0
rect 1030 -1200 1080 0
rect 1130 -1200 1180 0
rect 1360 -1200 1410 0
rect 1460 -1200 1510 0
<< pmos >>
rect -270 1440 -220 2640
rect -70 1440 -20 2640
rect 30 1440 80 2640
rect 130 1440 180 2640
rect 230 1440 280 2640
rect 330 1440 380 2640
rect 430 1440 480 2640
rect 530 1440 580 2640
rect 630 1440 680 2640
rect 730 1440 780 2640
rect 830 1440 880 2640
rect 930 1440 980 2640
rect 1030 1440 1080 2640
rect 1130 1440 1180 2640
rect 1230 1440 1280 2640
rect 1430 1440 1480 2640
rect -300 -2500 -250 -1300
rect -200 -2500 -150 -1300
rect 30 -2500 80 -1300
rect 130 -2500 180 -1300
rect 230 -2500 280 -1300
rect 330 -2500 380 -1300
rect 430 -2500 480 -1300
rect 530 -2500 580 -1300
rect 630 -2500 680 -1300
rect 730 -2500 780 -1300
rect 830 -2500 880 -1300
rect 930 -2500 980 -1300
rect 1030 -2500 1080 -1300
rect 1130 -2500 1180 -1300
rect 1360 -2500 1410 -1300
rect 1460 -2500 1510 -1300
<< ndiff >>
rect -350 1325 -300 1340
rect -350 155 -335 1325
rect -315 155 -300 1325
rect -350 140 -300 155
rect -250 1325 -200 1340
rect -250 155 -235 1325
rect -215 155 -200 1325
rect -250 140 -200 155
rect -150 1325 -100 1340
rect -150 155 -135 1325
rect -115 155 -100 1325
rect -150 140 -100 155
rect -20 1325 30 1340
rect -20 155 -5 1325
rect 15 155 30 1325
rect -20 140 30 155
rect 80 1325 130 1340
rect 80 155 95 1325
rect 115 155 130 1325
rect 80 140 130 155
rect 180 140 230 1340
rect 280 140 330 1340
rect 380 140 430 1340
rect 480 140 530 1340
rect 580 1325 630 1340
rect 580 155 595 1325
rect 615 155 630 1325
rect 580 140 630 155
rect 680 140 730 1340
rect 780 140 830 1340
rect 880 140 930 1340
rect 980 140 1030 1340
rect 1080 1325 1130 1340
rect 1080 155 1095 1325
rect 1115 155 1130 1325
rect 1080 140 1130 155
rect 1180 1325 1230 1340
rect 1180 155 1195 1325
rect 1215 155 1230 1325
rect 1180 140 1230 155
rect 1310 1325 1360 1340
rect 1310 155 1325 1325
rect 1345 155 1360 1325
rect 1310 140 1360 155
rect 1410 1325 1460 1340
rect 1410 155 1425 1325
rect 1445 155 1460 1325
rect 1410 140 1460 155
rect 1510 1325 1560 1340
rect 1510 155 1525 1325
rect 1545 155 1560 1325
rect 1510 140 1560 155
rect -350 -15 -300 0
rect -350 -1185 -335 -15
rect -315 -1185 -300 -15
rect -350 -1200 -300 -1185
rect -250 -15 -200 0
rect -250 -1185 -235 -15
rect -215 -1185 -200 -15
rect -250 -1200 -200 -1185
rect -150 -15 -100 0
rect -150 -1185 -135 -15
rect -115 -1185 -100 -15
rect -150 -1200 -100 -1185
rect -20 -15 30 0
rect -20 -1185 -5 -15
rect 15 -1185 30 -15
rect -20 -1200 30 -1185
rect 80 -15 130 0
rect 80 -1185 95 -15
rect 115 -1185 130 -15
rect 80 -1200 130 -1185
rect 180 -15 230 0
rect 180 -1185 195 -15
rect 215 -1185 230 -15
rect 180 -1200 230 -1185
rect 280 -15 330 0
rect 280 -1185 295 -15
rect 315 -1185 330 -15
rect 280 -1200 330 -1185
rect 380 -15 430 0
rect 380 -1185 395 -15
rect 415 -1185 430 -15
rect 380 -1200 430 -1185
rect 480 -15 530 0
rect 480 -1185 495 -15
rect 515 -1185 530 -15
rect 480 -1200 530 -1185
rect 580 -15 630 0
rect 580 -1185 595 -15
rect 615 -1185 630 -15
rect 580 -1200 630 -1185
rect 680 -15 730 0
rect 680 -1185 695 -15
rect 715 -1185 730 -15
rect 680 -1200 730 -1185
rect 780 -15 830 0
rect 780 -1185 795 -15
rect 815 -1185 830 -15
rect 780 -1200 830 -1185
rect 880 -15 930 0
rect 880 -1185 895 -15
rect 915 -1185 930 -15
rect 880 -1200 930 -1185
rect 980 -15 1030 0
rect 980 -1185 995 -15
rect 1015 -1185 1030 -15
rect 980 -1200 1030 -1185
rect 1080 -15 1130 0
rect 1080 -1185 1095 -15
rect 1115 -1185 1130 -15
rect 1080 -1200 1130 -1185
rect 1180 -15 1230 0
rect 1180 -1185 1195 -15
rect 1215 -1185 1230 -15
rect 1180 -1200 1230 -1185
rect 1310 -15 1360 0
rect 1310 -1185 1325 -15
rect 1345 -1185 1360 -15
rect 1310 -1200 1360 -1185
rect 1410 -15 1460 0
rect 1410 -1185 1425 -15
rect 1445 -1185 1460 -15
rect 1410 -1200 1460 -1185
rect 1510 -15 1560 0
rect 1510 -1185 1525 -15
rect 1545 -1185 1560 -15
rect 1510 -1200 1560 -1185
<< pdiff >>
rect -320 2625 -270 2640
rect -320 1455 -305 2625
rect -285 1455 -270 2625
rect -320 1440 -270 1455
rect -220 2625 -170 2640
rect -120 2625 -70 2640
rect -220 1455 -205 2625
rect -185 1455 -170 2625
rect -120 1455 -105 2625
rect -85 1455 -70 2625
rect -220 1440 -170 1455
rect -120 1440 -70 1455
rect -20 2625 30 2640
rect -20 1455 -5 2625
rect 15 1455 30 2625
rect -20 1440 30 1455
rect 80 2625 130 2640
rect 80 1455 95 2625
rect 115 1455 130 2625
rect 80 1440 130 1455
rect 180 2625 230 2640
rect 180 1455 195 2625
rect 215 1455 230 2625
rect 180 1440 230 1455
rect 280 2625 330 2640
rect 280 1455 295 2625
rect 315 1455 330 2625
rect 280 1440 330 1455
rect 380 2625 430 2640
rect 380 1455 395 2625
rect 415 1455 430 2625
rect 380 1440 430 1455
rect 480 2625 530 2640
rect 480 1455 495 2625
rect 515 1455 530 2625
rect 480 1440 530 1455
rect 580 2625 630 2640
rect 580 1455 595 2625
rect 615 1455 630 2625
rect 580 1440 630 1455
rect 680 2625 730 2640
rect 680 1455 695 2625
rect 715 1455 730 2625
rect 680 1440 730 1455
rect 780 2625 830 2640
rect 780 1455 795 2625
rect 815 1455 830 2625
rect 780 1440 830 1455
rect 880 2625 930 2640
rect 880 1455 895 2625
rect 915 1455 930 2625
rect 880 1440 930 1455
rect 980 2625 1030 2640
rect 980 1455 995 2625
rect 1015 1455 1030 2625
rect 980 1440 1030 1455
rect 1080 2625 1130 2640
rect 1080 1455 1095 2625
rect 1115 1455 1130 2625
rect 1080 1440 1130 1455
rect 1180 2625 1230 2640
rect 1180 1455 1195 2625
rect 1215 1455 1230 2625
rect 1180 1440 1230 1455
rect 1280 2625 1330 2640
rect 1380 2625 1430 2640
rect 1280 1455 1295 2625
rect 1315 1455 1330 2625
rect 1380 1455 1395 2625
rect 1415 1455 1430 2625
rect 1280 1440 1330 1455
rect 1380 1440 1430 1455
rect 1480 2625 1530 2640
rect 1480 1455 1495 2625
rect 1515 1455 1530 2625
rect 1480 1440 1530 1455
rect -350 -1315 -300 -1300
rect -350 -2485 -335 -1315
rect -315 -2485 -300 -1315
rect -350 -2500 -300 -2485
rect -250 -1315 -200 -1300
rect -250 -2485 -235 -1315
rect -215 -2485 -200 -1315
rect -250 -2500 -200 -2485
rect -150 -1315 -100 -1300
rect -150 -2485 -135 -1315
rect -115 -2485 -100 -1315
rect -150 -2500 -100 -2485
rect -20 -1315 30 -1300
rect -20 -2485 -5 -1315
rect 15 -2485 30 -1315
rect -20 -2500 30 -2485
rect 80 -1315 130 -1300
rect 80 -2485 95 -1315
rect 115 -2485 130 -1315
rect 80 -2500 130 -2485
rect 180 -2500 230 -1300
rect 280 -2500 330 -1300
rect 380 -2500 430 -1300
rect 480 -2500 530 -1300
rect 580 -1315 630 -1300
rect 580 -2485 595 -1315
rect 615 -2485 630 -1315
rect 580 -2500 630 -2485
rect 680 -2500 730 -1300
rect 780 -2500 830 -1300
rect 880 -2500 930 -1300
rect 980 -2500 1030 -1300
rect 1080 -1315 1130 -1300
rect 1080 -2485 1095 -1315
rect 1115 -2485 1130 -1315
rect 1080 -2500 1130 -2485
rect 1180 -1315 1230 -1300
rect 1180 -2485 1195 -1315
rect 1215 -2485 1230 -1315
rect 1180 -2500 1230 -2485
rect 1310 -1315 1360 -1300
rect 1310 -2485 1325 -1315
rect 1345 -2485 1360 -1315
rect 1310 -2500 1360 -2485
rect 1410 -1315 1460 -1300
rect 1410 -2485 1425 -1315
rect 1445 -2485 1460 -1315
rect 1410 -2500 1460 -2485
rect 1510 -1315 1560 -1300
rect 1510 -2485 1525 -1315
rect 1545 -2485 1560 -1315
rect 1510 -2500 1560 -2485
<< ndiffc >>
rect -335 155 -315 1325
rect -235 155 -215 1325
rect -135 155 -115 1325
rect -5 155 15 1325
rect 95 155 115 1325
rect 595 155 615 1325
rect 1095 155 1115 1325
rect 1195 155 1215 1325
rect 1325 155 1345 1325
rect 1425 155 1445 1325
rect 1525 155 1545 1325
rect -335 -1185 -315 -15
rect -235 -1185 -215 -15
rect -135 -1185 -115 -15
rect -5 -1185 15 -15
rect 95 -1185 115 -15
rect 195 -1185 215 -15
rect 295 -1185 315 -15
rect 395 -1185 415 -15
rect 495 -1185 515 -15
rect 595 -1185 615 -15
rect 695 -1185 715 -15
rect 795 -1185 815 -15
rect 895 -1185 915 -15
rect 995 -1185 1015 -15
rect 1095 -1185 1115 -15
rect 1195 -1185 1215 -15
rect 1325 -1185 1345 -15
rect 1425 -1185 1445 -15
rect 1525 -1185 1545 -15
<< pdiffc >>
rect -305 1455 -285 2625
rect -205 1455 -185 2625
rect -105 1455 -85 2625
rect -5 1455 15 2625
rect 95 1455 115 2625
rect 195 1455 215 2625
rect 295 1455 315 2625
rect 395 1455 415 2625
rect 495 1455 515 2625
rect 595 1455 615 2625
rect 695 1455 715 2625
rect 795 1455 815 2625
rect 895 1455 915 2625
rect 995 1455 1015 2625
rect 1095 1455 1115 2625
rect 1195 1455 1215 2625
rect 1295 1455 1315 2625
rect 1395 1455 1415 2625
rect 1495 1455 1515 2625
rect -335 -2485 -315 -1315
rect -235 -2485 -215 -1315
rect -135 -2485 -115 -1315
rect -5 -2485 15 -1315
rect 95 -2485 115 -1315
rect 595 -2485 615 -1315
rect 1095 -2485 1115 -1315
rect 1195 -2485 1215 -1315
rect 1325 -2485 1345 -1315
rect 1425 -2485 1445 -1315
rect 1525 -2485 1545 -1315
<< psubdiff >>
rect -100 1325 -50 1340
rect -100 155 -85 1325
rect -65 155 -50 1325
rect -100 140 -50 155
rect 1260 1325 1310 1340
rect 1260 155 1275 1325
rect 1295 155 1310 1325
rect 1260 140 1310 155
rect -100 -15 -50 0
rect -100 -1185 -85 -15
rect -65 -1185 -50 -15
rect -100 -1200 -50 -1185
rect 1260 -15 1310 0
rect 1260 -1185 1275 -15
rect 1295 -1185 1310 -15
rect 1260 -1200 1310 -1185
<< nsubdiff >>
rect -170 2625 -120 2640
rect -170 1455 -155 2625
rect -135 1455 -120 2625
rect -170 1440 -120 1455
rect 1330 2625 1380 2640
rect 1330 1455 1345 2625
rect 1365 1455 1380 2625
rect 1330 1440 1380 1455
rect -100 -1315 -50 -1300
rect -100 -2485 -85 -1315
rect -65 -2485 -50 -1315
rect -100 -2500 -50 -2485
rect 1260 -1315 1310 -1300
rect 1260 -2485 1275 -1315
rect 1295 -2485 1310 -1315
rect 1260 -2500 1310 -2485
<< psubdiffcont >>
rect -85 155 -65 1325
rect 1275 155 1295 1325
rect -85 -1185 -65 -15
rect 1275 -1185 1295 -15
<< nsubdiffcont >>
rect -155 1455 -135 2625
rect 1345 1455 1365 2625
rect -85 -2485 -65 -1315
rect 1275 -2485 1295 -1315
<< poly >>
rect -270 2640 -220 2655
rect -70 2640 -20 2655
rect 30 2640 80 2655
rect 130 2640 180 2655
rect 230 2640 280 2655
rect 330 2640 380 2655
rect 430 2640 480 2655
rect 530 2640 580 2655
rect 630 2640 680 2655
rect 730 2640 780 2655
rect 830 2640 880 2655
rect 930 2640 980 2655
rect 1030 2640 1080 2655
rect 1130 2640 1180 2655
rect 1230 2640 1280 2655
rect 1430 2640 1480 2655
rect -270 1425 -220 1440
rect -70 1425 -20 1440
rect -270 1415 -170 1425
rect -270 1405 -205 1415
rect -350 1385 -300 1400
rect -350 1365 -335 1385
rect -315 1375 -300 1385
rect -220 1395 -205 1405
rect -185 1395 -170 1415
rect -220 1380 -170 1395
rect -120 1415 -20 1425
rect -120 1395 -105 1415
rect -85 1405 -20 1415
rect 30 1415 80 1440
rect -85 1395 -70 1405
rect -120 1380 -70 1395
rect 30 1395 45 1415
rect 65 1395 80 1415
rect 30 1385 80 1395
rect 130 1415 180 1440
rect 130 1395 145 1415
rect 165 1395 180 1415
rect 130 1385 180 1395
rect 230 1415 280 1440
rect 230 1395 245 1415
rect 265 1395 280 1415
rect 230 1385 280 1395
rect 330 1415 380 1440
rect 330 1395 345 1415
rect 365 1395 380 1415
rect 330 1385 380 1395
rect 430 1415 480 1440
rect 430 1395 445 1415
rect 465 1395 480 1415
rect 430 1385 480 1395
rect 530 1415 580 1440
rect 530 1395 545 1415
rect 565 1395 580 1415
rect 530 1385 580 1395
rect 630 1415 680 1440
rect 630 1395 645 1415
rect 665 1395 680 1415
rect 630 1385 680 1395
rect 730 1415 780 1440
rect 730 1395 745 1415
rect 765 1395 780 1415
rect 730 1385 780 1395
rect 830 1415 880 1440
rect 830 1395 845 1415
rect 865 1395 880 1415
rect 830 1385 880 1395
rect 930 1415 980 1440
rect 930 1395 945 1415
rect 965 1395 980 1415
rect 930 1385 980 1395
rect 1030 1415 1080 1440
rect 1030 1395 1045 1415
rect 1065 1395 1080 1415
rect 1030 1385 1080 1395
rect 1130 1415 1180 1440
rect 1130 1395 1145 1415
rect 1165 1395 1180 1415
rect 1230 1425 1280 1440
rect 1430 1425 1480 1440
rect 1230 1415 1325 1425
rect 1230 1405 1290 1415
rect 1130 1385 1180 1395
rect 1275 1395 1290 1405
rect 1310 1395 1325 1415
rect 1275 1380 1325 1395
rect 1380 1415 1480 1425
rect 1380 1395 1395 1415
rect 1415 1410 1480 1415
rect 1415 1395 1430 1410
rect 1380 1380 1430 1395
rect 1510 1385 1560 1400
rect -315 1365 -250 1375
rect 1510 1370 1525 1385
rect -350 1355 -250 1365
rect 1460 1365 1525 1370
rect 1545 1365 1560 1385
rect 1460 1355 1560 1365
rect -300 1340 -250 1355
rect -200 1340 -150 1355
rect 30 1340 80 1355
rect 130 1340 180 1355
rect 230 1340 280 1355
rect 330 1340 380 1355
rect 430 1340 480 1355
rect 530 1340 580 1355
rect 630 1340 680 1355
rect 730 1340 780 1355
rect 830 1340 880 1355
rect 930 1340 980 1355
rect 1030 1340 1080 1355
rect 1130 1340 1180 1355
rect 1360 1340 1410 1355
rect 1460 1340 1510 1355
rect -300 120 -250 140
rect -200 95 -150 140
rect 30 120 80 140
rect 130 120 180 140
rect 230 120 280 140
rect 330 120 380 140
rect 430 120 480 140
rect 530 120 580 140
rect 630 120 680 140
rect 730 120 780 140
rect 830 120 880 140
rect 930 120 980 140
rect 1030 120 1080 140
rect 1130 120 1180 140
rect 30 100 1180 120
rect 30 95 80 100
rect -200 85 80 95
rect -200 65 -185 85
rect -165 80 80 85
rect 1130 95 1180 100
rect 1360 95 1410 140
rect 1460 120 1510 140
rect 1130 85 1580 95
rect 1130 80 1375 85
rect -165 65 -150 80
rect -300 0 -250 15
rect -200 0 -150 65
rect 1360 65 1375 80
rect 1395 80 1580 85
rect 1395 65 1410 80
rect 30 0 80 15
rect 130 0 180 15
rect 230 0 280 15
rect 330 0 380 15
rect 430 0 480 15
rect 530 0 580 15
rect 630 0 680 15
rect 730 0 780 15
rect 830 0 880 15
rect 930 0 980 15
rect 1030 0 1080 15
rect 1130 0 1180 15
rect 1360 0 1410 65
rect 1510 40 1560 55
rect 1510 35 1525 40
rect 1460 20 1525 35
rect 1545 20 1560 40
rect 1460 10 1560 20
rect 1460 0 1510 10
rect -300 -1215 -250 -1200
rect -200 -1215 -150 -1200
rect -350 -1225 -250 -1215
rect -350 -1245 -335 -1225
rect -315 -1235 -250 -1225
rect 30 -1225 80 -1200
rect -315 -1245 -300 -1235
rect -350 -1260 -300 -1245
rect 30 -1245 45 -1225
rect 65 -1245 80 -1225
rect 30 -1260 80 -1245
rect 130 -1225 180 -1200
rect 130 -1245 145 -1225
rect 165 -1245 180 -1225
rect 130 -1260 180 -1245
rect 230 -1225 280 -1200
rect 230 -1245 245 -1225
rect 265 -1245 280 -1225
rect 230 -1260 280 -1245
rect 330 -1225 380 -1200
rect 330 -1245 345 -1225
rect 365 -1245 380 -1225
rect 330 -1260 380 -1245
rect 430 -1225 480 -1200
rect 430 -1245 445 -1225
rect 465 -1245 480 -1225
rect 430 -1260 480 -1245
rect 530 -1225 580 -1200
rect 530 -1245 545 -1225
rect 565 -1245 580 -1225
rect 530 -1260 580 -1245
rect 630 -1225 680 -1200
rect 630 -1245 645 -1225
rect 665 -1245 680 -1225
rect 630 -1260 680 -1245
rect 730 -1225 780 -1200
rect 730 -1245 745 -1225
rect 765 -1245 780 -1225
rect 730 -1260 780 -1245
rect 830 -1225 880 -1200
rect 830 -1245 845 -1225
rect 865 -1245 880 -1225
rect 830 -1260 880 -1245
rect 930 -1225 980 -1200
rect 930 -1245 945 -1225
rect 965 -1245 980 -1225
rect 930 -1260 980 -1245
rect 1030 -1225 1080 -1200
rect 1030 -1245 1045 -1225
rect 1065 -1245 1080 -1225
rect 1030 -1260 1080 -1245
rect 1130 -1225 1180 -1200
rect 1360 -1215 1410 -1200
rect 1460 -1215 1510 -1200
rect 1130 -1245 1145 -1225
rect 1165 -1245 1180 -1225
rect 1130 -1260 1580 -1245
rect -300 -1300 -250 -1285
rect -200 -1300 -150 -1285
rect 30 -1300 80 -1285
rect 130 -1300 180 -1285
rect 230 -1300 280 -1285
rect 330 -1300 380 -1285
rect 430 -1300 480 -1285
rect 530 -1300 580 -1285
rect 630 -1300 680 -1285
rect 730 -1300 780 -1285
rect 830 -1300 880 -1285
rect 930 -1300 980 -1285
rect 1030 -1300 1080 -1285
rect 1130 -1300 1180 -1285
rect 1360 -1300 1410 -1285
rect 1460 -1300 1510 -1285
rect -300 -2515 -250 -2500
rect -350 -2525 -250 -2515
rect -350 -2545 -335 -2525
rect -315 -2535 -250 -2525
rect -200 -2515 -150 -2500
rect 30 -2515 80 -2500
rect 130 -2515 180 -2500
rect 230 -2515 280 -2500
rect 330 -2515 380 -2500
rect 430 -2515 480 -2500
rect 530 -2515 580 -2500
rect 630 -2515 680 -2500
rect 730 -2515 780 -2500
rect 830 -2515 880 -2500
rect 930 -2515 980 -2500
rect 1030 -2515 1080 -2500
rect 1130 -2515 1180 -2500
rect 1360 -2515 1410 -2500
rect -200 -2525 1410 -2515
rect -315 -2545 -300 -2535
rect -350 -2560 -300 -2545
rect -200 -2545 -185 -2525
rect -165 -2530 1375 -2525
rect -165 -2545 -150 -2530
rect -200 -2560 -150 -2545
rect 1360 -2545 1375 -2530
rect 1395 -2545 1410 -2525
rect 1460 -2515 1510 -2500
rect 1460 -2525 1560 -2515
rect 1460 -2535 1525 -2525
rect 1360 -2560 1410 -2545
rect 1510 -2545 1525 -2535
rect 1545 -2545 1560 -2525
rect 1510 -2560 1560 -2545
<< polycont >>
rect -335 1365 -315 1385
rect -205 1395 -185 1415
rect -105 1395 -85 1415
rect 45 1395 65 1415
rect 145 1395 165 1415
rect 245 1395 265 1415
rect 345 1395 365 1415
rect 445 1395 465 1415
rect 545 1395 565 1415
rect 645 1395 665 1415
rect 745 1395 765 1415
rect 845 1395 865 1415
rect 945 1395 965 1415
rect 1045 1395 1065 1415
rect 1145 1395 1165 1415
rect 1290 1395 1310 1415
rect 1395 1395 1415 1415
rect 1525 1365 1545 1385
rect -185 65 -165 85
rect 1375 65 1395 85
rect 1525 20 1545 40
rect -335 -1245 -315 -1225
rect 45 -1245 65 -1225
rect 145 -1245 165 -1225
rect 245 -1245 265 -1225
rect 345 -1245 365 -1225
rect 445 -1245 465 -1225
rect 545 -1245 565 -1225
rect 645 -1245 665 -1225
rect 745 -1245 765 -1225
rect 845 -1245 865 -1225
rect 945 -1245 965 -1225
rect 1045 -1245 1065 -1225
rect 1145 -1245 1165 -1225
rect -335 -2545 -315 -2525
rect -185 -2545 -165 -2525
rect 1375 -2545 1395 -2525
rect 1525 -2545 1545 -2525
<< locali >>
rect -315 2655 25 2675
rect -315 2625 -275 2655
rect -315 1455 -305 2625
rect -285 1455 -275 2625
rect -315 1445 -275 1455
rect -215 2625 -75 2635
rect -215 1455 -205 2625
rect -185 1455 -155 2625
rect -135 1455 -105 2625
rect -85 1455 -75 2625
rect -215 1445 -75 1455
rect -215 1425 -175 1445
rect -115 1425 -75 1445
rect -15 2625 25 2655
rect -15 1455 -5 2625
rect 15 1455 25 2625
rect -15 1425 25 1455
rect 85 2655 525 2675
rect 85 2625 125 2655
rect 85 1455 95 2625
rect 115 1455 125 2625
rect 85 1445 125 1455
rect 185 2625 225 2635
rect 185 1455 195 2625
rect 215 1455 225 2625
rect 185 1425 225 1455
rect 285 2625 325 2655
rect 285 1455 295 2625
rect 315 1455 325 2625
rect 285 1445 325 1455
rect 385 2625 425 2635
rect 385 1455 395 2625
rect 415 1455 425 2625
rect 385 1425 425 1455
rect 485 2625 525 2655
rect 685 2655 1125 2675
rect 485 1455 495 2625
rect 515 1455 525 2625
rect 485 1445 525 1455
rect 585 2625 625 2635
rect 585 1455 595 2625
rect 615 1455 625 2625
rect 585 1445 625 1455
rect 685 2625 725 2655
rect 685 1455 695 2625
rect 715 1455 725 2625
rect 685 1445 725 1455
rect 785 2625 825 2635
rect 785 1455 795 2625
rect 815 1455 825 2625
rect 785 1425 825 1455
rect 885 2625 925 2655
rect 885 1455 895 2625
rect 915 1455 925 2625
rect 885 1445 925 1455
rect 985 2625 1025 2635
rect 985 1455 995 2625
rect 1015 1455 1025 2625
rect 985 1425 1025 1455
rect 1085 2625 1125 2655
rect 1085 1455 1095 2625
rect 1115 1455 1125 2625
rect 1085 1445 1125 1455
rect 1185 2655 1525 2675
rect 1185 2625 1225 2655
rect 1185 1455 1195 2625
rect 1215 1455 1225 2625
rect 1185 1425 1225 1455
rect 1285 2625 1425 2635
rect 1285 1455 1295 2625
rect 1315 1455 1345 2625
rect 1365 1455 1395 2625
rect 1415 1455 1425 2625
rect 1285 1445 1425 1455
rect 1485 2625 1525 2655
rect 1485 1455 1495 2625
rect 1515 1455 1525 2625
rect 1485 1445 1525 1455
rect 1285 1425 1325 1445
rect 1385 1425 1425 1445
rect -220 1415 -170 1425
rect -220 1395 -205 1415
rect -185 1395 -170 1415
rect -350 1385 -300 1395
rect -220 1385 -170 1395
rect -120 1415 -70 1425
rect -120 1395 -105 1415
rect -85 1395 -70 1415
rect -120 1385 -70 1395
rect -15 1415 80 1425
rect -15 1395 45 1415
rect 65 1395 80 1415
rect -15 1385 80 1395
rect 130 1415 1080 1425
rect 130 1395 145 1415
rect 165 1395 245 1415
rect 265 1395 345 1415
rect 365 1395 445 1415
rect 465 1395 545 1415
rect 565 1395 645 1415
rect 665 1395 745 1415
rect 765 1395 845 1415
rect 865 1395 945 1415
rect 965 1395 1045 1415
rect 1065 1395 1080 1415
rect 130 1385 1080 1395
rect 1130 1415 1225 1425
rect 1130 1395 1145 1415
rect 1165 1395 1225 1415
rect 1130 1385 1225 1395
rect 1275 1415 1325 1425
rect 1275 1395 1290 1415
rect 1310 1395 1325 1415
rect 1275 1385 1325 1395
rect 1380 1415 1430 1425
rect 1380 1395 1395 1415
rect 1415 1395 1430 1415
rect 1380 1385 1430 1395
rect 1510 1385 1560 1395
rect -350 1365 -335 1385
rect -315 1365 -300 1385
rect -350 1355 -300 1365
rect -345 1325 -305 1355
rect -345 155 -335 1325
rect -315 155 -305 1325
rect -345 145 -305 155
rect -245 1325 -205 1335
rect -245 155 -235 1325
rect -215 155 -205 1325
rect -245 95 -205 155
rect -145 1325 -55 1335
rect -145 155 -135 1325
rect -115 155 -85 1325
rect -65 155 -55 1325
rect -145 145 -55 155
rect -15 1325 25 1385
rect -15 155 -5 1325
rect 15 155 25 1325
rect -15 145 25 155
rect 85 1325 125 1335
rect 85 155 95 1325
rect 115 155 125 1325
rect 85 145 125 155
rect 585 1325 625 1385
rect 585 155 595 1325
rect 615 155 625 1325
rect 585 145 625 155
rect 1085 1325 1125 1335
rect 1085 155 1095 1325
rect 1115 155 1125 1325
rect 1085 145 1125 155
rect 1185 1325 1225 1385
rect 1510 1365 1525 1385
rect 1545 1365 1560 1385
rect 1510 1355 1560 1365
rect 1185 155 1195 1325
rect 1215 155 1225 1325
rect -245 85 -150 95
rect -245 65 -185 85
rect -165 65 -150 85
rect -245 55 -150 65
rect 1185 35 1225 155
rect 1265 1325 1355 1335
rect 1265 155 1275 1325
rect 1295 155 1325 1325
rect 1345 155 1355 1325
rect 1265 145 1355 155
rect 1415 1325 1455 1335
rect 1415 155 1425 1325
rect 1445 155 1455 1325
rect 1415 145 1455 155
rect 1515 1325 1555 1355
rect 1515 155 1525 1325
rect 1545 155 1555 1325
rect 1515 145 1555 155
rect 1415 95 1445 145
rect 1360 85 1445 95
rect 1360 65 1375 85
rect 1395 65 1445 85
rect 1360 55 1445 65
rect 1470 70 1580 90
rect 1470 35 1490 70
rect 85 15 525 35
rect -345 -15 -305 -5
rect -345 -1185 -335 -15
rect -315 -1185 -305 -15
rect -345 -1215 -305 -1185
rect -245 -15 -205 -5
rect -245 -1185 -235 -15
rect -215 -1185 -205 -15
rect -350 -1225 -300 -1215
rect -350 -1245 -335 -1225
rect -315 -1245 -300 -1225
rect -350 -1255 -300 -1245
rect -345 -1315 -305 -1305
rect -345 -2485 -335 -1315
rect -315 -2485 -305 -1315
rect -345 -2515 -305 -2485
rect -245 -1315 -205 -1185
rect -145 -15 -55 -5
rect -145 -1185 -135 -15
rect -115 -1185 -85 -15
rect -65 -1185 -55 -15
rect -145 -1195 -55 -1185
rect -15 -15 25 -5
rect -15 -1185 -5 -15
rect 15 -1185 25 -15
rect -15 -1215 25 -1185
rect 85 -15 125 15
rect 85 -1185 95 -15
rect 115 -1185 125 -15
rect 85 -1195 125 -1185
rect 185 -15 225 -5
rect 185 -1185 195 -15
rect 215 -1185 225 -15
rect 185 -1215 225 -1185
rect 285 -15 325 15
rect 285 -1185 295 -15
rect 315 -1185 325 -15
rect 285 -1195 325 -1185
rect 385 -15 425 -5
rect 385 -1185 395 -15
rect 415 -1185 425 -15
rect 385 -1215 425 -1185
rect 485 -15 525 15
rect 685 15 1125 35
rect 1185 15 1490 35
rect 1510 40 1560 50
rect 1510 20 1525 40
rect 1545 20 1560 40
rect 485 -1185 495 -15
rect 515 -1185 525 -15
rect 485 -1195 525 -1185
rect 585 -15 625 -5
rect 585 -1185 595 -15
rect 615 -1185 625 -15
rect 585 -1195 625 -1185
rect 685 -15 725 15
rect 685 -1185 695 -15
rect 715 -1185 725 -15
rect 685 -1195 725 -1185
rect 785 -15 825 -5
rect 785 -1185 795 -15
rect 815 -1185 825 -15
rect 785 -1215 825 -1185
rect 885 -15 925 15
rect 885 -1185 895 -15
rect 915 -1185 925 -15
rect 885 -1195 925 -1185
rect 985 -15 1025 -5
rect 985 -1185 995 -15
rect 1015 -1185 1025 -15
rect 985 -1215 1025 -1185
rect 1085 -15 1125 15
rect 1510 10 1560 20
rect 1085 -1185 1095 -15
rect 1115 -1185 1125 -15
rect 1085 -1195 1125 -1185
rect 1185 -15 1225 -5
rect 1185 -1185 1195 -15
rect 1215 -1185 1225 -15
rect 1185 -1215 1225 -1185
rect 1265 -15 1355 -5
rect 1265 -1185 1275 -15
rect 1295 -1185 1325 -15
rect 1345 -1185 1355 -15
rect 1265 -1195 1355 -1185
rect 1415 -15 1455 -5
rect 1415 -1185 1425 -15
rect 1445 -1185 1455 -15
rect -15 -1225 80 -1215
rect -15 -1245 45 -1225
rect 65 -1245 80 -1225
rect -15 -1255 80 -1245
rect 130 -1225 1080 -1215
rect 130 -1245 145 -1225
rect 165 -1245 245 -1225
rect 265 -1245 345 -1225
rect 365 -1245 445 -1225
rect 465 -1245 545 -1225
rect 565 -1245 645 -1225
rect 665 -1245 745 -1225
rect 765 -1245 845 -1225
rect 865 -1245 945 -1225
rect 965 -1245 1045 -1225
rect 1065 -1245 1080 -1225
rect 130 -1255 1080 -1245
rect 1130 -1225 1225 -1215
rect 1130 -1245 1145 -1225
rect 1165 -1245 1225 -1225
rect 1130 -1255 1225 -1245
rect -245 -2485 -235 -1315
rect -215 -2485 -205 -1315
rect -245 -2515 -205 -2485
rect -145 -1315 -55 -1305
rect -145 -2485 -135 -1315
rect -115 -2485 -85 -1315
rect -65 -2485 -55 -1315
rect -145 -2495 -55 -2485
rect -15 -1315 25 -1255
rect -15 -2485 -5 -1315
rect 15 -2485 25 -1315
rect -15 -2495 25 -2485
rect 85 -1315 125 -1305
rect 85 -2485 95 -1315
rect 115 -2485 125 -1315
rect 85 -2495 125 -2485
rect 585 -1315 625 -1255
rect 585 -2485 595 -1315
rect 615 -2485 625 -1315
rect 585 -2495 625 -2485
rect 1085 -1315 1125 -1305
rect 1085 -2485 1095 -1315
rect 1115 -2485 1125 -1315
rect 1085 -2495 1125 -2485
rect 1185 -1315 1225 -1255
rect 1415 -1255 1455 -1185
rect 1515 -15 1555 10
rect 1515 -1185 1525 -15
rect 1545 -1185 1555 -15
rect 1515 -1195 1555 -1185
rect 1415 -1275 1580 -1255
rect 1185 -2485 1195 -1315
rect 1215 -2485 1225 -1315
rect 1185 -2495 1225 -2485
rect 1265 -1315 1355 -1305
rect 1265 -2485 1275 -1315
rect 1295 -2485 1325 -1315
rect 1345 -2485 1355 -1315
rect 1265 -2495 1355 -2485
rect 1415 -1315 1455 -1275
rect 1415 -2485 1425 -1315
rect 1445 -2485 1455 -1315
rect 1415 -2515 1455 -2485
rect 1515 -1315 1555 -1305
rect 1515 -2485 1525 -1315
rect 1545 -2485 1555 -1315
rect 1515 -2515 1555 -2485
rect -350 -2525 -300 -2515
rect -350 -2545 -335 -2525
rect -315 -2545 -300 -2525
rect -350 -2555 -300 -2545
rect -245 -2525 -150 -2515
rect -245 -2545 -185 -2525
rect -165 -2545 -150 -2525
rect -245 -2555 -150 -2545
rect 1360 -2525 1455 -2515
rect 1360 -2545 1375 -2525
rect 1395 -2545 1455 -2525
rect 1360 -2555 1455 -2545
rect 1510 -2525 1560 -2515
rect 1510 -2545 1525 -2525
rect 1545 -2545 1560 -2525
rect 1510 -2555 1560 -2545
<< viali >>
rect -205 1455 -185 2625
rect -155 1455 -135 2625
rect -105 1455 -85 2625
rect 595 1455 615 2625
rect 1295 1455 1315 2625
rect 1345 1455 1365 2625
rect 1395 1455 1415 2625
rect -335 155 -315 1325
rect -135 155 -115 1325
rect -85 155 -65 1325
rect 95 155 115 1325
rect 1095 155 1115 1325
rect 1275 155 1295 1325
rect 1325 155 1345 1325
rect 1525 155 1545 1325
rect -335 -1185 -315 -15
rect -335 -2485 -315 -1315
rect -135 -1185 -115 -15
rect -85 -1185 -65 -15
rect 595 -1185 615 -15
rect 1275 -1185 1295 -15
rect 1325 -1185 1345 -15
rect -135 -2485 -115 -1315
rect -85 -2485 -65 -1315
rect 95 -2485 115 -1315
rect 1095 -2485 1115 -1315
rect 1525 -1185 1545 -15
rect 1275 -2485 1295 -1315
rect 1325 -2485 1345 -1315
rect 1525 -2485 1545 -1315
<< metal1 >>
rect -370 2625 1580 2635
rect -370 1455 -205 2625
rect -185 1455 -155 2625
rect -135 1455 -105 2625
rect -85 1455 595 2625
rect 615 1455 1295 2625
rect 1315 1455 1345 2625
rect 1365 1455 1395 2625
rect 1415 1455 1580 2625
rect -370 1445 1580 1455
rect 1460 1335 1560 1340
rect -370 1325 1580 1335
rect -370 155 -335 1325
rect -315 155 -135 1325
rect -115 155 -85 1325
rect -65 155 95 1325
rect 115 155 1095 1325
rect 1115 155 1275 1325
rect 1295 155 1325 1325
rect 1345 155 1525 1325
rect 1545 155 1580 1325
rect -370 -15 1580 155
rect -370 -1185 -335 -15
rect -315 -1185 -135 -15
rect -115 -1185 -85 -15
rect -65 -1185 595 -15
rect 615 -1185 1275 -15
rect 1295 -1185 1325 -15
rect 1345 -1185 1525 -15
rect 1545 -1185 1580 -15
rect -370 -1195 1580 -1185
rect -370 -1315 1580 -1305
rect -370 -2485 -335 -1315
rect -315 -2485 -135 -1315
rect -115 -2485 -85 -1315
rect -65 -2485 95 -1315
rect 115 -2485 1095 -1315
rect 1115 -2485 1275 -1315
rect 1295 -2485 1325 -1315
rect 1345 -2485 1525 -1315
rect 1545 -2485 1580 -1315
rect -370 -2495 1580 -2485
<< labels >>
rlabel metal1 -370 2050 -370 2050 7 VP
port 6 w
rlabel locali 1580 80 1580 80 3 Vcp
port 3 e
rlabel locali 1580 -1265 1580 -1265 3 Vbp
port 5 e
rlabel poly 1580 -1250 1580 -1250 3 Vcn
port 10 e
rlabel metal1 -370 -1900 -370 -1900 7 VP
port 9 w
rlabel metal1 -370 50 -370 50 7 VN
port 7 w
rlabel poly 1580 90 1580 90 3 Vbn
port 8 e
<< end >>
