magic
tech sky130A
timestamp 1697774992
<< nwell >>
rect -270 1420 1480 2670
rect -270 -2485 1480 -1245
<< nmos >>
rect -200 145 -150 1345
rect 30 145 80 1345
rect 130 145 180 1345
rect 230 145 280 1345
rect 330 145 380 1345
rect 430 145 480 1345
rect 530 145 580 1345
rect 630 145 680 1345
rect 730 145 780 1345
rect 830 145 880 1345
rect 930 145 980 1345
rect 1030 145 1080 1345
rect 1130 145 1180 1345
rect 1360 145 1410 1345
rect -200 -1165 -150 35
rect 30 -1165 80 35
rect 130 -1165 180 35
rect 230 -1165 280 35
rect 330 -1165 380 35
rect 430 -1165 480 35
rect 530 -1165 580 35
rect 630 -1165 680 35
rect 730 -1165 780 35
rect 830 -1165 880 35
rect 930 -1165 980 35
rect 1030 -1165 1080 35
rect 1130 -1165 1180 35
rect 1360 -1165 1410 35
<< pmos >>
rect -70 1440 -20 2640
rect 30 1440 80 2640
rect 130 1440 180 2640
rect 230 1440 280 2640
rect 330 1440 380 2640
rect 430 1440 480 2640
rect 530 1440 580 2640
rect 630 1440 680 2640
rect 730 1440 780 2640
rect 830 1440 880 2640
rect 930 1440 980 2640
rect 1030 1440 1080 2640
rect 1130 1440 1180 2640
rect 1230 1440 1280 2640
rect -200 -2465 -150 -1265
rect 30 -2465 80 -1265
rect 130 -2465 180 -1265
rect 230 -2465 280 -1265
rect 330 -2465 380 -1265
rect 430 -2465 480 -1265
rect 530 -2465 580 -1265
rect 630 -2465 680 -1265
rect 730 -2465 780 -1265
rect 830 -2465 880 -1265
rect 930 -2465 980 -1265
rect 1030 -2465 1080 -1265
rect 1130 -2465 1180 -1265
rect 1360 -2465 1410 -1265
<< ndiff >>
rect -250 1330 -200 1345
rect -250 160 -235 1330
rect -215 160 -200 1330
rect -250 145 -200 160
rect -150 1330 -100 1345
rect -150 160 -135 1330
rect -115 160 -100 1330
rect -150 145 -100 160
rect -20 1330 30 1345
rect -20 160 -5 1330
rect 15 160 30 1330
rect -20 145 30 160
rect 80 1330 130 1345
rect 80 160 95 1330
rect 115 160 130 1330
rect 80 145 130 160
rect 180 145 230 1345
rect 280 145 330 1345
rect 380 145 430 1345
rect 480 145 530 1345
rect 580 1330 630 1345
rect 580 160 595 1330
rect 615 160 630 1330
rect 580 145 630 160
rect 680 145 730 1345
rect 780 145 830 1345
rect 880 145 930 1345
rect 980 145 1030 1345
rect 1080 1330 1130 1345
rect 1080 160 1095 1330
rect 1115 160 1130 1330
rect 1080 145 1130 160
rect 1180 1330 1230 1345
rect 1180 160 1195 1330
rect 1215 160 1230 1330
rect 1180 145 1230 160
rect 1310 1330 1360 1345
rect 1310 160 1325 1330
rect 1345 160 1360 1330
rect 1310 145 1360 160
rect 1410 1330 1460 1345
rect 1410 160 1425 1330
rect 1445 160 1460 1330
rect 1410 145 1460 160
rect -250 20 -200 35
rect -250 -1150 -235 20
rect -215 -1150 -200 20
rect -250 -1165 -200 -1150
rect -150 20 -100 35
rect -150 -1150 -135 20
rect -115 -1150 -100 20
rect -150 -1165 -100 -1150
rect -20 20 30 35
rect -20 -1150 -5 20
rect 15 -1150 30 20
rect -20 -1165 30 -1150
rect 80 20 130 35
rect 80 -1150 95 20
rect 115 -1150 130 20
rect 80 -1165 130 -1150
rect 180 20 230 35
rect 180 -1150 195 20
rect 215 -1150 230 20
rect 180 -1165 230 -1150
rect 280 20 330 35
rect 280 -1150 295 20
rect 315 -1150 330 20
rect 280 -1165 330 -1150
rect 380 20 430 35
rect 380 -1150 395 20
rect 415 -1150 430 20
rect 380 -1165 430 -1150
rect 480 20 530 35
rect 480 -1150 495 20
rect 515 -1150 530 20
rect 480 -1165 530 -1150
rect 580 20 630 35
rect 580 -1150 595 20
rect 615 -1150 630 20
rect 580 -1165 630 -1150
rect 680 20 730 35
rect 680 -1150 695 20
rect 715 -1150 730 20
rect 680 -1165 730 -1150
rect 780 20 830 35
rect 780 -1150 795 20
rect 815 -1150 830 20
rect 780 -1165 830 -1150
rect 880 20 930 35
rect 880 -1150 895 20
rect 915 -1150 930 20
rect 880 -1165 930 -1150
rect 980 20 1030 35
rect 980 -1150 995 20
rect 1015 -1150 1030 20
rect 980 -1165 1030 -1150
rect 1080 20 1130 35
rect 1080 -1150 1095 20
rect 1115 -1150 1130 20
rect 1080 -1165 1130 -1150
rect 1180 20 1230 35
rect 1180 -1150 1195 20
rect 1215 -1150 1230 20
rect 1180 -1165 1230 -1150
rect 1310 20 1360 35
rect 1310 -1150 1325 20
rect 1345 -1150 1360 20
rect 1310 -1165 1360 -1150
rect 1410 20 1460 35
rect 1410 -1150 1425 20
rect 1445 -1150 1460 20
rect 1410 -1165 1460 -1150
<< pdiff >>
rect -120 2625 -70 2640
rect -120 1455 -105 2625
rect -85 1455 -70 2625
rect -120 1440 -70 1455
rect -20 2625 30 2640
rect -20 1455 -5 2625
rect 15 1455 30 2625
rect -20 1440 30 1455
rect 80 2625 130 2640
rect 80 1455 95 2625
rect 115 1455 130 2625
rect 80 1440 130 1455
rect 180 2625 230 2640
rect 180 1455 195 2625
rect 215 1455 230 2625
rect 180 1440 230 1455
rect 280 2625 330 2640
rect 280 1455 295 2625
rect 315 1455 330 2625
rect 280 1440 330 1455
rect 380 2625 430 2640
rect 380 1455 395 2625
rect 415 1455 430 2625
rect 380 1440 430 1455
rect 480 2625 530 2640
rect 480 1455 495 2625
rect 515 1455 530 2625
rect 480 1440 530 1455
rect 580 2625 630 2640
rect 580 1455 595 2625
rect 615 1455 630 2625
rect 580 1440 630 1455
rect 680 2625 730 2640
rect 680 1455 695 2625
rect 715 1455 730 2625
rect 680 1440 730 1455
rect 780 2625 830 2640
rect 780 1455 795 2625
rect 815 1455 830 2625
rect 780 1440 830 1455
rect 880 2625 930 2640
rect 880 1455 895 2625
rect 915 1455 930 2625
rect 880 1440 930 1455
rect 980 2625 1030 2640
rect 980 1455 995 2625
rect 1015 1455 1030 2625
rect 980 1440 1030 1455
rect 1080 2625 1130 2640
rect 1080 1455 1095 2625
rect 1115 1455 1130 2625
rect 1080 1440 1130 1455
rect 1180 2625 1230 2640
rect 1180 1455 1195 2625
rect 1215 1455 1230 2625
rect 1180 1440 1230 1455
rect 1280 2625 1330 2640
rect 1280 1455 1295 2625
rect 1315 1455 1330 2625
rect 1280 1440 1330 1455
rect -250 -1280 -200 -1265
rect -250 -2450 -235 -1280
rect -215 -2450 -200 -1280
rect -250 -2465 -200 -2450
rect -150 -1280 -100 -1265
rect -150 -2450 -135 -1280
rect -115 -2450 -100 -1280
rect -150 -2465 -100 -2450
rect -20 -1280 30 -1265
rect -20 -2450 -5 -1280
rect 15 -2450 30 -1280
rect -20 -2465 30 -2450
rect 80 -1280 130 -1265
rect 80 -2450 95 -1280
rect 115 -2450 130 -1280
rect 80 -2465 130 -2450
rect 180 -2465 230 -1265
rect 280 -2465 330 -1265
rect 380 -2465 430 -1265
rect 480 -2465 530 -1265
rect 580 -1280 630 -1265
rect 580 -2450 595 -1280
rect 615 -2450 630 -1280
rect 580 -2465 630 -2450
rect 680 -2465 730 -1265
rect 780 -2465 830 -1265
rect 880 -2465 930 -1265
rect 980 -2465 1030 -1265
rect 1080 -1280 1130 -1265
rect 1080 -2450 1095 -1280
rect 1115 -2450 1130 -1280
rect 1080 -2465 1130 -2450
rect 1180 -1280 1230 -1265
rect 1180 -2450 1195 -1280
rect 1215 -2450 1230 -1280
rect 1180 -2465 1230 -2450
rect 1310 -1280 1360 -1265
rect 1310 -2450 1325 -1280
rect 1345 -2450 1360 -1280
rect 1310 -2465 1360 -2450
rect 1410 -1280 1460 -1265
rect 1410 -2450 1425 -1280
rect 1445 -2450 1460 -1280
rect 1410 -2465 1460 -2450
<< ndiffc >>
rect -235 160 -215 1330
rect -135 160 -115 1330
rect -5 160 15 1330
rect 95 160 115 1330
rect 595 160 615 1330
rect 1095 160 1115 1330
rect 1195 160 1215 1330
rect 1325 160 1345 1330
rect 1425 160 1445 1330
rect -235 -1150 -215 20
rect -135 -1150 -115 20
rect -5 -1150 15 20
rect 95 -1150 115 20
rect 195 -1150 215 20
rect 295 -1150 315 20
rect 395 -1150 415 20
rect 495 -1150 515 20
rect 595 -1150 615 20
rect 695 -1150 715 20
rect 795 -1150 815 20
rect 895 -1150 915 20
rect 995 -1150 1015 20
rect 1095 -1150 1115 20
rect 1195 -1150 1215 20
rect 1325 -1150 1345 20
rect 1425 -1150 1445 20
<< pdiffc >>
rect -105 1455 -85 2625
rect -5 1455 15 2625
rect 95 1455 115 2625
rect 195 1455 215 2625
rect 295 1455 315 2625
rect 395 1455 415 2625
rect 495 1455 515 2625
rect 595 1455 615 2625
rect 695 1455 715 2625
rect 795 1455 815 2625
rect 895 1455 915 2625
rect 995 1455 1015 2625
rect 1095 1455 1115 2625
rect 1195 1455 1215 2625
rect 1295 1455 1315 2625
rect -235 -2450 -215 -1280
rect -135 -2450 -115 -1280
rect -5 -2450 15 -1280
rect 95 -2450 115 -1280
rect 595 -2450 615 -1280
rect 1095 -2450 1115 -1280
rect 1195 -2450 1215 -1280
rect 1325 -2450 1345 -1280
rect 1425 -2450 1445 -1280
<< psubdiff >>
rect -100 1330 -50 1345
rect -100 160 -85 1330
rect -65 160 -50 1330
rect -100 145 -50 160
rect 1260 1330 1310 1345
rect 1260 160 1275 1330
rect 1295 160 1310 1330
rect 1260 145 1310 160
rect -100 20 -50 35
rect -100 -1150 -85 20
rect -65 -1150 -50 20
rect -100 -1165 -50 -1150
rect 1260 20 1310 35
rect 1260 -1150 1275 20
rect 1295 -1150 1310 20
rect 1260 -1165 1310 -1150
<< nsubdiff >>
rect -170 2625 -120 2640
rect -170 1455 -155 2625
rect -135 1455 -120 2625
rect -170 1440 -120 1455
rect 1330 2625 1380 2640
rect 1330 1455 1345 2625
rect 1365 1455 1380 2625
rect 1330 1440 1380 1455
rect -100 -1280 -50 -1265
rect -100 -2450 -85 -1280
rect -65 -2450 -50 -1280
rect -100 -2465 -50 -2450
rect 1260 -1280 1310 -1265
rect 1260 -2450 1275 -1280
rect 1295 -2450 1310 -1280
rect 1260 -2465 1310 -2450
<< psubdiffcont >>
rect -85 160 -65 1330
rect 1275 160 1295 1330
rect -85 -1150 -65 20
rect 1275 -1150 1295 20
<< nsubdiffcont >>
rect -155 1455 -135 2625
rect 1345 1455 1365 2625
rect -85 -2450 -65 -1280
rect 1275 -2450 1295 -1280
<< poly >>
rect -70 2640 -20 2655
rect 30 2640 80 2655
rect 130 2640 180 2655
rect 230 2640 280 2655
rect 330 2640 380 2655
rect 430 2640 480 2655
rect 530 2640 580 2655
rect 630 2640 680 2655
rect 730 2640 780 2655
rect 830 2640 880 2655
rect 930 2640 980 2655
rect 1030 2640 1080 2655
rect 1130 2640 1180 2655
rect 1230 2640 1280 2655
rect -70 1425 -20 1440
rect -120 1415 -20 1425
rect -120 1395 -105 1415
rect -85 1405 -20 1415
rect 30 1415 80 1440
rect -85 1395 -70 1405
rect -120 1380 -70 1395
rect 30 1395 45 1415
rect 65 1395 80 1415
rect 30 1385 80 1395
rect 130 1415 180 1440
rect 130 1395 145 1415
rect 165 1395 180 1415
rect 130 1385 180 1395
rect 230 1415 280 1440
rect 230 1395 245 1415
rect 265 1395 280 1415
rect 230 1385 280 1395
rect 330 1415 380 1440
rect 330 1395 345 1415
rect 365 1395 380 1415
rect 330 1385 380 1395
rect 430 1415 480 1440
rect 430 1395 445 1415
rect 465 1395 480 1415
rect 430 1385 480 1395
rect 530 1415 580 1440
rect 530 1395 545 1415
rect 565 1395 580 1415
rect 530 1385 580 1395
rect 630 1415 680 1440
rect 630 1395 645 1415
rect 665 1395 680 1415
rect 630 1385 680 1395
rect 730 1415 780 1440
rect 730 1395 745 1415
rect 765 1395 780 1415
rect 730 1385 780 1395
rect 830 1415 880 1440
rect 830 1395 845 1415
rect 865 1395 880 1415
rect 830 1385 880 1395
rect 930 1415 980 1440
rect 930 1395 945 1415
rect 965 1395 980 1415
rect 930 1385 980 1395
rect 1030 1415 1080 1440
rect 1030 1395 1045 1415
rect 1065 1395 1080 1415
rect 1030 1385 1080 1395
rect 1130 1415 1180 1440
rect 1130 1395 1145 1415
rect 1165 1395 1180 1415
rect 1230 1425 1280 1440
rect 1230 1415 1325 1425
rect 1230 1405 1290 1415
rect 1130 1385 1180 1395
rect 1275 1395 1290 1405
rect 1310 1395 1325 1415
rect 1275 1380 1325 1395
rect -200 1345 -150 1360
rect 30 1345 80 1360
rect 130 1345 180 1360
rect 230 1345 280 1360
rect 330 1345 380 1360
rect 430 1345 480 1360
rect 530 1345 580 1360
rect 630 1345 680 1360
rect 730 1345 780 1360
rect 830 1345 880 1360
rect 930 1345 980 1360
rect 1030 1345 1080 1360
rect 1130 1345 1180 1360
rect 1360 1345 1410 1360
rect -200 130 -150 145
rect 30 130 80 145
rect 130 130 180 145
rect 230 130 280 145
rect 330 130 380 145
rect 430 130 480 145
rect 530 130 580 145
rect 630 130 680 145
rect 730 130 780 145
rect 830 130 880 145
rect 930 130 980 145
rect 1030 130 1080 145
rect 1130 130 1180 145
rect 1360 130 1410 145
rect -200 120 1480 130
rect -200 100 -185 120
rect -165 115 1375 120
rect -165 100 -150 115
rect -200 35 -150 100
rect 1360 100 1375 115
rect 1395 115 1480 120
rect 1395 100 1410 115
rect 30 35 80 50
rect 130 35 180 50
rect 230 35 280 50
rect 330 35 380 50
rect 430 35 480 50
rect 530 35 580 50
rect 630 35 680 50
rect 730 35 780 50
rect 830 35 880 50
rect 930 35 980 50
rect 1030 35 1080 50
rect 1130 35 1180 50
rect 1360 35 1410 100
rect -200 -1180 -150 -1165
rect 30 -1190 80 -1165
rect 30 -1210 45 -1190
rect 65 -1210 80 -1190
rect 30 -1225 80 -1210
rect 130 -1190 180 -1165
rect 130 -1210 145 -1190
rect 165 -1210 180 -1190
rect 130 -1225 180 -1210
rect 230 -1190 280 -1165
rect 230 -1210 245 -1190
rect 265 -1210 280 -1190
rect 230 -1225 280 -1210
rect 330 -1190 380 -1165
rect 330 -1210 345 -1190
rect 365 -1210 380 -1190
rect 330 -1225 380 -1210
rect 430 -1190 480 -1165
rect 430 -1210 445 -1190
rect 465 -1210 480 -1190
rect 430 -1225 480 -1210
rect 530 -1190 580 -1165
rect 530 -1210 545 -1190
rect 565 -1210 580 -1190
rect 530 -1225 580 -1210
rect 630 -1190 680 -1165
rect 630 -1210 645 -1190
rect 665 -1210 680 -1190
rect 630 -1225 680 -1210
rect 730 -1190 780 -1165
rect 730 -1210 745 -1190
rect 765 -1210 780 -1190
rect 730 -1225 780 -1210
rect 830 -1190 880 -1165
rect 830 -1210 845 -1190
rect 865 -1210 880 -1190
rect 830 -1225 880 -1210
rect 930 -1190 980 -1165
rect 930 -1210 945 -1190
rect 965 -1210 980 -1190
rect 930 -1225 980 -1210
rect 1030 -1190 1080 -1165
rect 1030 -1210 1045 -1190
rect 1065 -1210 1080 -1190
rect 1030 -1225 1080 -1210
rect 1130 -1190 1180 -1165
rect 1360 -1180 1410 -1165
rect 1130 -1210 1145 -1190
rect 1165 -1210 1180 -1190
rect 1130 -1225 1480 -1210
rect -200 -1265 -150 -1250
rect 30 -1265 80 -1250
rect 130 -1265 180 -1250
rect 230 -1265 280 -1250
rect 330 -1265 380 -1250
rect 430 -1265 480 -1250
rect 530 -1265 580 -1250
rect 630 -1265 680 -1250
rect 730 -1265 780 -1250
rect 830 -1265 880 -1250
rect 930 -1265 980 -1250
rect 1030 -1265 1080 -1250
rect 1130 -1265 1180 -1250
rect 1360 -1265 1410 -1250
rect -200 -2480 -150 -2465
rect 30 -2480 80 -2465
rect 130 -2480 180 -2465
rect 230 -2480 280 -2465
rect 330 -2480 380 -2465
rect 430 -2480 480 -2465
rect 530 -2480 580 -2465
rect 630 -2480 680 -2465
rect 730 -2480 780 -2465
rect 830 -2480 880 -2465
rect 930 -2480 980 -2465
rect 1030 -2480 1080 -2465
rect 1130 -2480 1180 -2465
rect 1360 -2480 1410 -2465
rect -200 -2490 1410 -2480
rect -200 -2510 -185 -2490
rect -165 -2495 1410 -2490
rect -165 -2510 -150 -2495
rect -200 -2525 -150 -2510
rect 1360 -2505 1410 -2495
rect 1360 -2525 1375 -2505
rect 1395 -2525 1410 -2505
rect 1360 -2540 1410 -2525
<< polycont >>
rect -105 1395 -85 1415
rect 45 1395 65 1415
rect 145 1395 165 1415
rect 245 1395 265 1415
rect 345 1395 365 1415
rect 445 1395 465 1415
rect 545 1395 565 1415
rect 645 1395 665 1415
rect 745 1395 765 1415
rect 845 1395 865 1415
rect 945 1395 965 1415
rect 1045 1395 1065 1415
rect 1145 1395 1165 1415
rect 1290 1395 1310 1415
rect -185 100 -165 120
rect 1375 100 1395 120
rect 45 -1210 65 -1190
rect 145 -1210 165 -1190
rect 245 -1210 265 -1190
rect 345 -1210 365 -1190
rect 445 -1210 465 -1190
rect 545 -1210 565 -1190
rect 645 -1210 665 -1190
rect 745 -1210 765 -1190
rect 845 -1210 865 -1190
rect 945 -1210 965 -1190
rect 1045 -1210 1065 -1190
rect 1145 -1210 1165 -1190
rect -185 -2510 -165 -2490
rect 1375 -2525 1395 -2505
<< locali >>
rect 85 2655 525 2675
rect -165 2625 -75 2635
rect -165 1455 -155 2625
rect -135 1455 -105 2625
rect -85 1455 -75 2625
rect -165 1445 -75 1455
rect -115 1425 -75 1445
rect -15 2625 25 2635
rect -15 1455 -5 2625
rect 15 1455 25 2625
rect -15 1425 25 1455
rect 85 2625 125 2655
rect 85 1455 95 2625
rect 115 1455 125 2625
rect 85 1445 125 1455
rect 185 2625 225 2635
rect 185 1455 195 2625
rect 215 1455 225 2625
rect 185 1425 225 1455
rect 285 2625 325 2655
rect 285 1455 295 2625
rect 315 1455 325 2625
rect 285 1445 325 1455
rect 385 2625 425 2635
rect 385 1455 395 2625
rect 415 1455 425 2625
rect 385 1425 425 1455
rect 485 2625 525 2655
rect 685 2655 1125 2675
rect 485 1455 495 2625
rect 515 1455 525 2625
rect 485 1445 525 1455
rect 585 2625 625 2635
rect 585 1455 595 2625
rect 615 1455 625 2625
rect 585 1445 625 1455
rect 685 2625 725 2655
rect 685 1455 695 2625
rect 715 1455 725 2625
rect 685 1445 725 1455
rect 785 2625 825 2635
rect 785 1455 795 2625
rect 815 1455 825 2625
rect 785 1425 825 1455
rect 885 2625 925 2655
rect 885 1455 895 2625
rect 915 1455 925 2625
rect 885 1445 925 1455
rect 985 2625 1025 2635
rect 985 1455 995 2625
rect 1015 1455 1025 2625
rect 985 1425 1025 1455
rect 1085 2625 1125 2655
rect 1085 1455 1095 2625
rect 1115 1455 1125 2625
rect 1085 1445 1125 1455
rect 1185 2625 1225 2635
rect 1185 1455 1195 2625
rect 1215 1455 1225 2625
rect 1185 1425 1225 1455
rect 1285 2625 1375 2635
rect 1285 1455 1295 2625
rect 1315 1455 1345 2625
rect 1365 1455 1375 2625
rect 1285 1445 1375 1455
rect 1285 1425 1325 1445
rect -120 1415 -70 1425
rect -120 1395 -105 1415
rect -85 1395 -70 1415
rect -120 1385 -70 1395
rect -15 1415 80 1425
rect -15 1395 45 1415
rect 65 1395 80 1415
rect -15 1385 80 1395
rect 130 1415 1080 1425
rect 130 1395 145 1415
rect 165 1395 245 1415
rect 265 1395 345 1415
rect 365 1395 445 1415
rect 465 1395 545 1415
rect 565 1395 645 1415
rect 665 1395 745 1415
rect 765 1395 845 1415
rect 865 1395 945 1415
rect 965 1395 1045 1415
rect 1065 1395 1080 1415
rect 130 1385 1080 1395
rect 1130 1415 1225 1425
rect 1130 1395 1145 1415
rect 1165 1395 1225 1415
rect 1130 1385 1225 1395
rect 1275 1415 1325 1425
rect 1275 1395 1290 1415
rect 1310 1395 1325 1415
rect 1275 1385 1325 1395
rect -245 1330 -205 1340
rect -245 160 -235 1330
rect -215 160 -205 1330
rect -245 130 -205 160
rect -145 1330 -55 1340
rect -145 160 -135 1330
rect -115 160 -85 1330
rect -65 160 -55 1330
rect -145 150 -55 160
rect -15 1330 25 1385
rect -15 160 -5 1330
rect 15 160 25 1330
rect -15 150 25 160
rect 85 1330 125 1340
rect 85 160 95 1330
rect 115 160 125 1330
rect 85 150 125 160
rect 585 1330 625 1385
rect 585 160 595 1330
rect 615 160 625 1330
rect 585 150 625 160
rect 1085 1330 1125 1340
rect 1085 160 1095 1330
rect 1115 160 1125 1330
rect 1085 150 1125 160
rect 1185 1330 1225 1385
rect 1185 160 1195 1330
rect 1215 160 1225 1330
rect -245 120 -150 130
rect -245 100 -185 120
rect -165 100 -150 120
rect -245 90 -150 100
rect 1185 70 1225 160
rect 1265 1330 1355 1340
rect 1265 160 1275 1330
rect 1295 160 1325 1330
rect 1345 160 1355 1330
rect 1265 150 1355 160
rect 1415 1330 1455 1340
rect 1415 160 1425 1330
rect 1445 160 1455 1330
rect 1415 130 1455 160
rect 1360 120 1455 130
rect 1360 100 1375 120
rect 1395 100 1455 120
rect 1360 90 1455 100
rect 85 50 525 70
rect -245 20 -205 30
rect -245 -1150 -235 20
rect -215 -1150 -205 20
rect -245 -1280 -205 -1150
rect -145 20 -55 30
rect -145 -1150 -135 20
rect -115 -1150 -85 20
rect -65 -1150 -55 20
rect -145 -1160 -55 -1150
rect -15 20 25 30
rect -15 -1150 -5 20
rect 15 -1150 25 20
rect -15 -1180 25 -1150
rect 85 20 125 50
rect 85 -1150 95 20
rect 115 -1150 125 20
rect 85 -1160 125 -1150
rect 185 20 225 30
rect 185 -1150 195 20
rect 215 -1150 225 20
rect 185 -1180 225 -1150
rect 285 20 325 50
rect 285 -1150 295 20
rect 315 -1150 325 20
rect 285 -1160 325 -1150
rect 385 20 425 30
rect 385 -1150 395 20
rect 415 -1150 425 20
rect 385 -1180 425 -1150
rect 485 20 525 50
rect 685 50 1125 70
rect 1185 50 1480 70
rect 485 -1150 495 20
rect 515 -1150 525 20
rect 485 -1160 525 -1150
rect 585 20 625 30
rect 585 -1150 595 20
rect 615 -1150 625 20
rect 585 -1160 625 -1150
rect 685 20 725 50
rect 685 -1150 695 20
rect 715 -1150 725 20
rect 685 -1160 725 -1150
rect 785 20 825 30
rect 785 -1150 795 20
rect 815 -1150 825 20
rect 785 -1180 825 -1150
rect 885 20 925 50
rect 885 -1150 895 20
rect 915 -1150 925 20
rect 885 -1160 925 -1150
rect 985 20 1025 30
rect 985 -1150 995 20
rect 1015 -1150 1025 20
rect 985 -1180 1025 -1150
rect 1085 20 1125 50
rect 1085 -1150 1095 20
rect 1115 -1150 1125 20
rect 1085 -1160 1125 -1150
rect 1185 20 1225 30
rect 1185 -1150 1195 20
rect 1215 -1150 1225 20
rect 1185 -1180 1225 -1150
rect 1265 20 1355 30
rect 1265 -1150 1275 20
rect 1295 -1150 1325 20
rect 1345 -1150 1355 20
rect 1265 -1160 1355 -1150
rect 1415 20 1455 30
rect 1415 -1150 1425 20
rect 1445 -1150 1455 20
rect -15 -1190 80 -1180
rect -15 -1210 45 -1190
rect 65 -1210 80 -1190
rect -15 -1220 80 -1210
rect 130 -1190 1080 -1180
rect 130 -1210 145 -1190
rect 165 -1210 245 -1190
rect 265 -1210 345 -1190
rect 365 -1210 445 -1190
rect 465 -1210 545 -1190
rect 565 -1210 645 -1190
rect 665 -1210 745 -1190
rect 765 -1210 845 -1190
rect 865 -1210 945 -1190
rect 965 -1210 1045 -1190
rect 1065 -1210 1080 -1190
rect 130 -1220 1080 -1210
rect 1130 -1190 1225 -1180
rect 1130 -1210 1145 -1190
rect 1165 -1210 1225 -1190
rect 1130 -1220 1225 -1210
rect -245 -2450 -235 -1280
rect -215 -2450 -205 -1280
rect -245 -2480 -205 -2450
rect -145 -1280 -55 -1270
rect -145 -2450 -135 -1280
rect -115 -2450 -85 -1280
rect -65 -2450 -55 -1280
rect -145 -2460 -55 -2450
rect -15 -1280 25 -1220
rect -15 -2450 -5 -1280
rect 15 -2450 25 -1280
rect -15 -2460 25 -2450
rect 85 -1280 125 -1270
rect 85 -2450 95 -1280
rect 115 -2450 125 -1280
rect 85 -2460 125 -2450
rect 585 -1280 625 -1220
rect 585 -2450 595 -1280
rect 615 -2450 625 -1280
rect 585 -2460 625 -2450
rect 1085 -1280 1125 -1270
rect 1085 -2450 1095 -1280
rect 1115 -2450 1125 -1280
rect 1085 -2460 1125 -2450
rect 1185 -1280 1225 -1220
rect 1415 -1220 1455 -1150
rect 1415 -1240 1480 -1220
rect 1185 -2450 1195 -1280
rect 1215 -2450 1225 -1280
rect 1185 -2460 1225 -2450
rect 1265 -1280 1355 -1270
rect 1265 -2450 1275 -1280
rect 1295 -2450 1325 -1280
rect 1345 -2450 1355 -1280
rect 1265 -2460 1355 -2450
rect 1415 -1280 1455 -1240
rect 1415 -2450 1425 -1280
rect 1445 -2450 1455 -1280
rect -245 -2490 -150 -2480
rect -245 -2510 -185 -2490
rect -165 -2510 -150 -2490
rect 1415 -2495 1455 -2450
rect -245 -2520 -150 -2510
rect 1360 -2505 1455 -2495
rect 1360 -2525 1375 -2505
rect 1395 -2525 1455 -2505
rect 1360 -2535 1455 -2525
<< viali >>
rect -155 1455 -135 2625
rect -105 1455 -85 2625
rect 595 1455 615 2625
rect 1295 1455 1315 2625
rect 1345 1455 1365 2625
rect -135 160 -115 1330
rect -85 160 -65 1330
rect 95 160 115 1330
rect 1095 160 1115 1330
rect 1275 160 1295 1330
rect 1325 160 1345 1330
rect -135 -1150 -115 20
rect -85 -1150 -65 20
rect 595 -1150 615 20
rect 1275 -1150 1295 20
rect 1325 -1150 1345 20
rect -135 -2450 -115 -1280
rect -85 -2450 -65 -1280
rect 95 -2450 115 -1280
rect 1095 -2450 1115 -1280
rect 1275 -2450 1295 -1280
rect 1325 -2450 1345 -1280
<< metal1 >>
rect -270 2625 1480 2635
rect -270 1455 -155 2625
rect -135 1455 -105 2625
rect -85 1455 595 2625
rect 615 1455 1295 2625
rect 1315 1455 1345 2625
rect 1365 1455 1480 2625
rect -270 1445 1480 1455
rect -270 1330 1480 1340
rect -270 160 -135 1330
rect -115 160 -85 1330
rect -65 160 95 1330
rect 115 160 1095 1330
rect 1115 160 1275 1330
rect 1295 160 1325 1330
rect 1345 160 1480 1330
rect -270 20 1480 160
rect -270 -1150 -135 20
rect -115 -1150 -85 20
rect -65 -1150 595 20
rect 615 -1150 1275 20
rect 1295 -1150 1325 20
rect 1345 -1150 1480 20
rect -270 -1160 1480 -1150
rect -270 -1280 1480 -1270
rect -270 -2450 -135 -1280
rect -115 -2450 -85 -1280
rect -65 -2450 95 -1280
rect 115 -2450 1095 -1280
rect 1115 -2450 1275 -1280
rect 1295 -2450 1325 -1280
rect 1345 -2450 1480 -1280
rect -270 -2460 1480 -2450
<< labels >>
rlabel metal1 -270 2050 -270 2050 7 VP
port 6 w
rlabel locali 1480 60 1480 60 3 Vcp
port 3 e
rlabel poly 1480 125 1480 125 3 Vbn
port 2 e
rlabel metal1 -270 -1865 -270 -1865 7 VP
port 9 w
rlabel locali 1480 -1230 1480 -1230 3 Vbp
port 5 e
rlabel poly 1480 -1215 1480 -1215 3 Vcn
port 10 e
rlabel metal1 -270 85 -270 85 7 VN
port 7 w
<< end >>
