magic
tech sky130A
timestamp 1695615073
<< nwell >>
rect -125 295 325 670
<< nmos >>
rect 70 100 85 200
rect 135 100 150 200
rect 200 100 215 200
rect -40 -135 -25 -35
rect 70 -135 85 -35
rect 135 -135 150 -35
rect 200 -135 215 -35
<< pmos >>
rect 0 550 15 650
rect 65 550 80 650
rect 130 550 145 650
rect 195 550 210 650
rect -50 315 -35 415
rect 15 315 30 415
rect 195 315 210 415
<< ndiff >>
rect 20 185 70 200
rect 20 115 35 185
rect 55 115 70 185
rect 20 100 70 115
rect 85 185 135 200
rect 85 115 100 185
rect 120 115 135 185
rect 85 100 135 115
rect 150 185 200 200
rect 150 115 165 185
rect 185 115 200 185
rect 150 100 200 115
rect 215 185 265 200
rect 215 115 230 185
rect 250 115 265 185
rect 215 100 265 115
rect -90 -50 -40 -35
rect -90 -120 -75 -50
rect -55 -120 -40 -50
rect -90 -135 -40 -120
rect -25 -50 70 -35
rect -25 -120 35 -50
rect 55 -120 70 -50
rect -25 -135 70 -120
rect 85 -50 135 -35
rect 85 -120 100 -50
rect 120 -120 135 -50
rect 85 -135 135 -120
rect 150 -50 200 -35
rect 150 -120 165 -50
rect 185 -120 200 -50
rect 150 -135 200 -120
rect 215 -50 265 -35
rect 215 -120 230 -50
rect 250 -120 265 -50
rect 215 -135 265 -120
<< pdiff >>
rect -50 635 0 650
rect -50 565 -35 635
rect -15 565 0 635
rect -50 550 0 565
rect 15 635 65 650
rect 15 565 30 635
rect 50 565 65 635
rect 15 550 65 565
rect 80 635 130 650
rect 80 565 95 635
rect 115 565 130 635
rect 80 550 130 565
rect 145 635 195 650
rect 145 565 160 635
rect 180 565 195 635
rect 145 550 195 565
rect 210 635 260 650
rect 210 565 225 635
rect 245 565 260 635
rect 210 550 260 565
rect -100 400 -50 415
rect -100 330 -85 400
rect -65 330 -50 400
rect -100 315 -50 330
rect -35 400 15 415
rect -35 330 -20 400
rect 0 330 15 400
rect -35 315 15 330
rect 30 400 80 415
rect 30 330 45 400
rect 65 330 80 400
rect 30 315 80 330
rect 145 400 195 415
rect 145 330 160 400
rect 180 330 195 400
rect 145 315 195 330
rect 210 400 260 415
rect 210 330 225 400
rect 245 330 260 400
rect 210 315 260 330
<< ndiffc >>
rect 35 115 55 185
rect 100 115 120 185
rect 165 115 185 185
rect 230 115 250 185
rect -75 -120 -55 -50
rect 35 -120 55 -50
rect 100 -120 120 -50
rect 165 -120 185 -50
rect 230 -120 250 -50
<< pdiffc >>
rect -35 565 -15 635
rect 30 565 50 635
rect 95 565 115 635
rect 160 565 180 635
rect 225 565 245 635
rect -85 330 -65 400
rect -20 330 0 400
rect 45 330 65 400
rect 160 330 180 400
rect 225 330 245 400
<< psubdiff >>
rect -30 185 20 200
rect -30 115 -15 185
rect 5 115 20 185
rect -30 100 20 115
<< nsubdiff >>
rect -100 635 -50 650
rect -100 565 -85 635
rect -65 565 -50 635
rect -100 550 -50 565
<< psubdiffcont >>
rect -15 115 5 185
<< nsubdiffcont >>
rect -85 565 -65 635
<< poly >>
rect 0 650 15 665
rect 65 650 80 665
rect 130 650 145 665
rect 195 650 210 665
rect 0 540 15 550
rect -50 525 15 540
rect -50 415 -35 525
rect 65 495 80 550
rect 130 535 145 550
rect 195 535 210 550
rect 195 525 235 535
rect 195 505 205 525
rect 225 505 235 525
rect 195 495 235 505
rect -10 485 80 495
rect -10 465 0 485
rect 20 480 80 485
rect 20 465 30 480
rect -10 455 30 465
rect 15 415 30 430
rect 195 415 210 430
rect -50 275 -35 315
rect -55 260 -35 275
rect 15 295 30 315
rect 15 285 55 295
rect 15 265 25 285
rect 45 270 55 285
rect 45 265 85 270
rect -55 80 -40 260
rect 15 255 85 265
rect 195 260 210 315
rect 70 200 85 255
rect 135 200 150 255
rect 195 250 235 260
rect 195 230 205 250
rect 225 230 235 250
rect 195 220 235 230
rect 200 200 215 220
rect 70 85 85 100
rect -55 65 -25 80
rect -40 -35 -25 65
rect 70 75 110 85
rect 70 55 80 75
rect 100 55 110 75
rect 70 45 110 55
rect 70 -35 85 45
rect 135 -35 150 100
rect 200 85 215 100
rect 200 50 240 60
rect 200 30 210 50
rect 230 30 240 50
rect 200 20 240 30
rect 200 -35 215 20
rect -40 -150 -25 -135
rect 70 -150 85 -135
rect 135 -150 150 -135
rect 200 -150 215 -135
<< polycont >>
rect 205 505 225 525
rect 0 465 20 485
rect 25 265 45 285
rect 205 230 225 250
rect 80 55 100 75
rect 210 30 230 50
<< locali >>
rect -95 635 -5 645
rect -95 565 -85 635
rect -65 565 -35 635
rect -15 565 -5 635
rect -95 555 -5 565
rect 20 635 60 645
rect 20 565 30 635
rect 50 565 60 635
rect 20 555 60 565
rect 85 635 125 645
rect 85 565 95 635
rect 115 565 125 635
rect 85 555 125 565
rect 150 635 190 645
rect 150 565 160 635
rect 180 565 190 635
rect 150 555 190 565
rect 215 635 255 645
rect 215 565 225 635
rect 245 575 255 635
rect 245 565 325 575
rect 215 555 325 565
rect -95 410 -75 555
rect 40 535 60 555
rect 40 515 115 535
rect -10 485 30 495
rect -10 465 0 485
rect 20 465 30 485
rect -10 455 30 465
rect -10 410 10 455
rect -95 400 -55 410
rect -95 330 -85 400
rect -65 330 -55 400
rect -95 320 -55 330
rect -30 400 10 410
rect -30 330 -20 400
rect 0 330 10 400
rect -30 320 10 330
rect 35 400 75 410
rect 35 330 45 400
rect 65 330 75 400
rect 35 320 75 330
rect 95 295 115 515
rect 195 525 235 535
rect 195 505 205 525
rect 225 505 235 525
rect 195 495 235 505
rect 215 410 235 495
rect 150 400 190 410
rect 150 330 160 400
rect 180 330 190 400
rect 150 320 190 330
rect 215 400 255 410
rect 215 330 225 400
rect 245 330 255 400
rect 215 320 255 330
rect 215 300 235 320
rect 15 285 115 295
rect 15 265 25 285
rect 45 275 115 285
rect 45 265 55 275
rect 15 255 55 265
rect 95 195 115 275
rect 155 280 235 300
rect 155 195 175 280
rect 280 260 300 555
rect 195 250 300 260
rect 195 230 205 250
rect 225 240 300 250
rect 225 230 235 240
rect 195 220 235 230
rect -25 185 65 195
rect -25 115 -15 185
rect 5 115 35 185
rect 55 115 65 185
rect -25 105 65 115
rect 90 185 130 195
rect 90 115 100 185
rect 120 115 130 185
rect 90 105 130 115
rect 155 185 195 195
rect 155 115 165 185
rect 185 115 195 185
rect 155 105 195 115
rect 220 185 260 195
rect 220 115 230 185
rect 250 115 260 185
rect 220 105 260 115
rect 25 -40 45 105
rect 90 85 110 105
rect 70 75 110 85
rect 70 55 80 75
rect 100 55 110 75
rect 70 45 110 55
rect 175 60 195 105
rect 175 50 240 60
rect 175 40 210 50
rect 200 30 210 40
rect 230 30 240 50
rect 200 20 240 30
rect 280 0 300 240
rect 175 -20 300 0
rect 175 -40 195 -20
rect -85 -50 -45 -40
rect -85 -120 -75 -50
rect -55 -120 -45 -50
rect -85 -130 -45 -120
rect 25 -50 65 -40
rect 25 -120 35 -50
rect 55 -120 65 -50
rect 25 -130 65 -120
rect 90 -50 130 -40
rect 90 -120 100 -50
rect 120 -120 130 -50
rect 90 -130 130 -120
rect 155 -50 195 -40
rect 155 -120 165 -50
rect 185 -120 195 -50
rect 155 -130 195 -120
rect 220 -50 260 -40
rect 220 -120 230 -50
rect 250 -120 260 -50
rect 220 -130 260 -120
<< end >>
