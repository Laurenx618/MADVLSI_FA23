magic
tech sky130A
timestamp 1695709979
<< nwell >>
rect -60 295 290 810
<< nmos >>
rect 10 -160 25 240
rect 75 140 90 240
rect 140 140 155 240
rect 205 140 220 240
rect 75 -125 90 -25
rect 140 -125 155 -25
rect 205 -125 220 -25
<< pmos >>
rect 10 615 25 715
rect 75 615 90 715
rect 10 315 25 415
rect 75 315 90 415
rect 150 315 165 715
rect 205 560 220 660
rect 205 315 220 415
<< ndiff >>
rect -40 225 10 240
rect -40 -145 -25 225
rect -5 -145 10 225
rect -40 -160 10 -145
rect 25 140 75 240
rect 90 225 140 240
rect 90 155 105 225
rect 125 155 140 225
rect 90 140 140 155
rect 155 225 205 240
rect 155 155 170 225
rect 190 155 205 225
rect 155 140 205 155
rect 220 225 270 240
rect 220 155 235 225
rect 255 155 270 225
rect 220 140 270 155
rect 25 -25 55 140
rect 25 -125 75 -25
rect 90 -40 140 -25
rect 90 -110 105 -40
rect 125 -110 140 -40
rect 90 -125 140 -110
rect 155 -40 205 -25
rect 155 -110 170 -40
rect 190 -110 205 -40
rect 155 -125 205 -110
rect 220 -40 270 -25
rect 220 -110 235 -40
rect 255 -110 270 -40
rect 220 -125 270 -110
rect 25 -160 55 -125
<< pdiff >>
rect -40 700 10 715
rect -40 630 -25 700
rect -5 630 10 700
rect -40 615 10 630
rect 25 700 75 715
rect 25 630 40 700
rect 60 630 75 700
rect 25 615 75 630
rect 90 700 150 715
rect 90 615 115 700
rect 100 415 115 615
rect -40 400 10 415
rect -40 330 -25 400
rect -5 330 10 400
rect -40 315 10 330
rect 25 400 75 415
rect 25 330 40 400
rect 60 330 75 400
rect 25 315 75 330
rect 90 330 115 415
rect 135 330 150 700
rect 90 315 150 330
rect 165 660 190 715
rect 165 560 205 660
rect 220 645 270 660
rect 220 575 235 645
rect 255 575 270 645
rect 220 560 270 575
rect 165 415 190 560
rect 165 315 205 415
rect 220 400 270 415
rect 220 330 235 400
rect 255 330 270 400
rect 220 315 270 330
<< ndiffc >>
rect -25 -145 -5 225
rect 105 155 125 225
rect 170 155 190 225
rect 235 155 255 225
rect 105 -110 125 -40
rect 170 -110 190 -40
rect 235 -110 255 -40
<< pdiffc >>
rect -25 630 -5 700
rect 40 630 60 700
rect -25 330 -5 400
rect 40 330 60 400
rect 115 330 135 700
rect 235 575 255 645
rect 235 330 255 400
<< psubdiff >>
rect 165 -170 280 -155
rect 165 -190 185 -170
rect 260 -190 280 -170
rect 165 -205 280 -190
<< nsubdiff >>
rect 220 770 270 790
rect 220 705 235 770
rect 255 705 270 770
rect 220 690 270 705
<< psubdiffcont >>
rect 185 -190 260 -170
<< nsubdiffcont >>
rect 235 705 255 770
<< poly >>
rect 10 755 165 770
rect 10 715 25 755
rect 75 715 90 730
rect 150 715 165 755
rect 10 605 25 615
rect 75 605 90 615
rect -60 590 25 605
rect 70 590 90 605
rect -60 440 -45 590
rect 70 560 85 590
rect -20 550 20 560
rect -20 530 -10 550
rect 10 530 20 550
rect -20 520 20 530
rect 45 550 85 560
rect 45 530 55 550
rect 75 530 85 550
rect 45 520 85 530
rect 5 480 20 520
rect 5 465 90 480
rect -60 425 25 440
rect 10 415 25 425
rect 75 415 90 465
rect 205 660 220 675
rect 205 545 220 560
rect 205 535 245 545
rect 205 515 215 535
rect 235 515 245 535
rect 205 505 245 515
rect 225 465 265 475
rect 225 450 235 465
rect 205 445 235 450
rect 255 445 265 465
rect 205 435 265 445
rect 205 415 220 435
rect 10 300 25 315
rect -15 290 25 300
rect -15 270 -5 290
rect 15 270 25 290
rect -15 260 25 270
rect 10 240 25 260
rect 75 240 90 315
rect 150 300 165 315
rect 140 285 165 300
rect 140 240 155 285
rect 205 240 220 315
rect 75 125 90 140
rect 75 115 115 125
rect 75 95 85 115
rect 105 95 115 115
rect 75 85 115 95
rect 65 50 105 60
rect 65 30 75 50
rect 95 30 105 50
rect 65 20 105 30
rect 75 -25 90 20
rect 140 -25 155 140
rect 205 125 220 140
rect 205 115 285 125
rect 205 110 255 115
rect 245 95 255 110
rect 275 95 285 115
rect 245 85 285 95
rect 180 75 220 85
rect 180 55 190 75
rect 210 55 220 75
rect 180 45 220 55
rect 205 -25 220 45
rect 75 -140 90 -125
rect 10 -175 25 -160
rect 140 -175 155 -125
rect 205 -140 220 -125
rect 10 -190 155 -175
<< polycont >>
rect -10 530 10 550
rect 55 530 75 550
rect 215 515 235 535
rect 235 445 255 465
rect -5 270 15 290
rect 85 95 105 115
rect 75 30 95 50
rect 255 95 275 115
rect 190 55 210 75
<< locali >>
rect 225 770 265 785
rect 225 750 235 770
rect 125 730 235 750
rect 125 710 145 730
rect -35 700 5 710
rect -35 640 -25 700
rect -60 630 -25 640
rect -5 630 5 700
rect -60 620 5 630
rect 30 700 70 710
rect 30 630 40 700
rect 60 630 70 700
rect 30 620 70 630
rect 105 700 145 710
rect 30 600 50 620
rect 0 580 50 600
rect 0 560 20 580
rect -20 550 20 560
rect -20 530 -10 550
rect 10 530 20 550
rect -20 520 20 530
rect 45 550 85 560
rect 45 530 55 550
rect 75 530 85 550
rect 45 520 85 530
rect 45 415 65 520
rect 45 410 70 415
rect -35 400 5 410
rect -35 340 -25 400
rect -60 330 -25 340
rect -5 330 5 400
rect -60 320 5 330
rect 30 400 70 410
rect 30 330 40 400
rect 60 330 70 400
rect 30 320 70 330
rect 105 330 115 700
rect 135 330 145 700
rect 225 705 235 730
rect 255 705 265 770
rect 225 695 265 705
rect 225 645 265 655
rect 225 575 235 645
rect 255 640 265 645
rect 255 620 290 640
rect 255 585 265 620
rect 255 575 285 585
rect 225 565 285 575
rect 205 535 245 545
rect 205 530 215 535
rect 105 320 145 330
rect 180 515 215 530
rect 235 515 245 535
rect 180 505 245 515
rect 180 410 200 505
rect 265 475 285 565
rect 225 465 285 475
rect 225 445 235 465
rect 255 455 285 465
rect 255 445 265 455
rect 225 435 265 445
rect 180 400 265 410
rect 180 390 235 400
rect -15 290 25 300
rect -15 280 -5 290
rect -60 270 -5 280
rect 15 270 25 290
rect -60 260 25 270
rect 50 235 70 320
rect 180 235 200 390
rect 225 330 235 390
rect 255 340 265 400
rect 255 330 290 340
rect 225 320 290 330
rect -35 225 5 235
rect -35 -145 -25 225
rect -5 -145 5 225
rect 35 225 135 235
rect 35 215 105 225
rect 35 60 55 215
rect 95 155 105 215
rect 125 155 135 225
rect 95 145 135 155
rect 160 225 200 235
rect 160 155 170 225
rect 190 155 200 225
rect 160 145 200 155
rect 225 225 265 235
rect 225 155 235 225
rect 255 155 265 225
rect 225 145 265 155
rect 75 115 115 125
rect 75 95 85 115
rect 105 105 115 115
rect 170 105 190 145
rect 245 115 285 125
rect 105 95 150 105
rect 75 85 150 95
rect 170 85 200 105
rect 245 95 255 115
rect 275 95 285 115
rect 245 85 285 95
rect 35 50 105 60
rect 35 40 75 50
rect 65 30 75 40
rect 95 30 105 50
rect 65 20 105 30
rect 130 5 150 85
rect 180 75 220 85
rect 180 55 190 75
rect 210 55 220 75
rect 180 45 220 55
rect 245 25 265 85
rect 115 -15 150 5
rect 180 5 265 25
rect 115 -30 135 -15
rect 180 -30 200 5
rect 95 -40 135 -30
rect 95 -110 105 -40
rect 125 -110 135 -40
rect 95 -120 135 -110
rect 160 -40 200 -30
rect 160 -110 170 -40
rect 190 -110 200 -40
rect 160 -120 200 -110
rect 225 -40 265 -30
rect 225 -110 235 -40
rect 255 -110 265 -40
rect 225 -120 265 -110
rect -35 -155 5 -145
rect 225 -160 245 -120
rect 170 -170 275 -160
rect 170 -190 185 -170
rect 260 -190 275 -170
rect 170 -200 275 -190
<< viali >>
rect 115 330 135 700
rect 235 705 255 770
rect -25 -145 -5 225
rect 235 -110 255 -40
rect 185 -190 260 -170
<< metal1 >>
rect -60 770 290 790
rect -60 705 235 770
rect 255 705 290 770
rect -60 700 290 705
rect -60 330 115 700
rect 135 330 290 700
rect -60 315 290 330
rect -60 225 290 240
rect -60 -145 -25 225
rect -5 -40 290 225
rect -5 -110 235 -40
rect 255 -110 290 -40
rect -5 -145 290 -110
rect -60 -170 290 -145
rect -60 -190 185 -170
rect 260 -190 290 -170
rect -60 -205 290 -190
<< labels >>
rlabel metal1 -60 30 -60 30 3 VN
port 7 e
rlabel locali -60 630 -60 630 7 D
port 1 w
rlabel locali -60 330 -60 330 7 DB
port 2 w
rlabel locali -60 270 -60 270 7 CLK
port 3 w
rlabel locali 290 630 290 630 3 Q
port 4 e
rlabel locali 290 330 290 330 3 QB
port 5 e
rlabel metal1 -60 560 -60 560 7 VP
port 6 w
<< end >>
