magic
tech sky130A
timestamp 1697676819
<< nwell >>
rect -730 1375 390 2625
<< nmos >>
rect -675 2695 -625 3895
rect -575 2695 -525 3895
rect -475 2695 -425 3895
rect -295 2695 -245 3895
rect -95 2695 -45 3895
rect 85 2695 135 3895
rect 185 2695 235 3895
rect 285 2695 335 3895
rect -625 15 -575 1215
rect -525 15 -475 1215
rect -425 15 -375 1215
rect -325 15 -275 1215
rect -65 15 -15 1215
rect 35 15 85 1215
rect 135 15 185 1215
rect 235 15 285 1215
<< pmos >>
rect -625 1400 -575 2600
rect -525 1400 -475 2600
rect -425 1400 -375 2600
rect -325 1400 -275 2600
rect -65 1400 -15 2600
rect 35 1400 85 2600
rect 135 1400 185 2600
rect 235 1400 285 2600
<< ndiff >>
rect -725 3880 -675 3895
rect -725 2710 -710 3880
rect -690 2710 -675 3880
rect -725 2695 -675 2710
rect -625 3880 -575 3895
rect -625 2710 -610 3880
rect -590 2710 -575 3880
rect -625 2695 -575 2710
rect -525 3880 -475 3895
rect -525 2710 -510 3880
rect -490 2710 -475 3880
rect -525 2695 -475 2710
rect -425 3880 -375 3895
rect -425 2710 -410 3880
rect -390 2710 -375 3880
rect -425 2695 -375 2710
rect -345 3880 -295 3895
rect -345 2710 -330 3880
rect -310 2710 -295 3880
rect -345 2695 -295 2710
rect -245 3880 -195 3895
rect -145 3880 -95 3895
rect -245 2710 -230 3880
rect -210 2710 -195 3880
rect -145 2710 -130 3880
rect -110 2710 -95 3880
rect -245 2695 -195 2710
rect -145 2695 -95 2710
rect -45 3880 5 3895
rect -45 2710 -30 3880
rect -10 2710 5 3880
rect -45 2695 5 2710
rect 35 3880 85 3895
rect 35 2710 50 3880
rect 70 2710 85 3880
rect 35 2695 85 2710
rect 135 3880 185 3895
rect 135 2710 150 3880
rect 170 2710 185 3880
rect 135 2695 185 2710
rect 235 3880 285 3895
rect 235 2710 250 3880
rect 270 2710 285 3880
rect 235 2695 285 2710
rect 335 3880 385 3895
rect 335 2710 350 3880
rect 370 2710 385 3880
rect 335 2695 385 2710
rect -675 1200 -625 1215
rect -675 30 -660 1200
rect -640 30 -625 1200
rect -675 15 -625 30
rect -575 15 -525 1215
rect -475 1200 -425 1215
rect -475 30 -460 1200
rect -440 30 -425 1200
rect -475 15 -425 30
rect -375 15 -325 1215
rect -275 1200 -225 1215
rect -275 30 -260 1200
rect -240 30 -225 1200
rect -275 15 -225 30
rect -115 1200 -65 1215
rect -115 30 -100 1200
rect -80 30 -65 1200
rect -115 15 -65 30
rect -15 15 35 1215
rect 85 1200 135 1215
rect 85 30 100 1200
rect 120 30 135 1200
rect 85 15 135 30
rect 185 15 235 1215
rect 285 1200 335 1215
rect 285 30 300 1200
rect 320 30 335 1200
rect 285 15 335 30
<< pdiff >>
rect -675 2585 -625 2600
rect -675 1415 -660 2585
rect -640 1415 -625 2585
rect -675 1400 -625 1415
rect -575 2585 -525 2600
rect -575 1415 -560 2585
rect -540 1415 -525 2585
rect -575 1400 -525 1415
rect -475 2585 -425 2600
rect -475 1415 -460 2585
rect -440 1415 -425 2585
rect -475 1400 -425 1415
rect -375 2585 -325 2600
rect -375 1415 -360 2585
rect -340 1415 -325 2585
rect -375 1400 -325 1415
rect -275 2585 -225 2600
rect -275 1415 -260 2585
rect -240 1415 -225 2585
rect -275 1400 -225 1415
rect -115 2585 -65 2600
rect -115 1415 -100 2585
rect -80 1415 -65 2585
rect -115 1400 -65 1415
rect -15 2585 35 2600
rect -15 1415 0 2585
rect 20 1415 35 2585
rect -15 1400 35 1415
rect 85 2585 135 2600
rect 85 1415 100 2585
rect 120 1415 135 2585
rect 85 1400 135 1415
rect 185 2585 235 2600
rect 185 1415 200 2585
rect 220 1415 235 2585
rect 185 1400 235 1415
rect 285 2585 335 2600
rect 285 1415 300 2585
rect 320 1415 335 2585
rect 285 1400 335 1415
<< ndiffc >>
rect -710 2710 -690 3880
rect -610 2710 -590 3880
rect -510 2710 -490 3880
rect -410 2710 -390 3880
rect -330 2710 -310 3880
rect -230 2710 -210 3880
rect -130 2710 -110 3880
rect -30 2710 -10 3880
rect 50 2710 70 3880
rect 150 2710 170 3880
rect 250 2710 270 3880
rect 350 2710 370 3880
rect -660 30 -640 1200
rect -460 30 -440 1200
rect -260 30 -240 1200
rect -100 30 -80 1200
rect 100 30 120 1200
rect 300 30 320 1200
<< pdiffc >>
rect -660 1415 -640 2585
rect -560 1415 -540 2585
rect -460 1415 -440 2585
rect -360 1415 -340 2585
rect -260 1415 -240 2585
rect -100 1415 -80 2585
rect 0 1415 20 2585
rect 100 1415 120 2585
rect 200 1415 220 2585
rect 300 1415 320 2585
<< psubdiff >>
rect -195 3880 -145 3895
rect -195 2710 -180 3880
rect -160 2710 -145 3880
rect -195 2695 -145 2710
rect -195 1200 -145 1215
rect -195 30 -180 1200
rect -160 30 -145 1200
rect -195 15 -145 30
<< nsubdiff >>
rect -195 2585 -145 2600
rect -195 1415 -180 2585
rect -160 1415 -145 2585
rect -195 1400 -145 1415
<< psubdiffcont >>
rect -180 2710 -160 3880
rect -180 30 -160 1200
<< nsubdiffcont >>
rect -180 1415 -160 2585
<< poly >>
rect -575 4025 390 4040
rect -725 3940 -675 3955
rect -725 3920 -710 3940
rect -690 3925 -675 3940
rect -690 3920 -625 3925
rect -725 3910 -625 3920
rect -675 3895 -625 3910
rect -575 3895 -525 4025
rect -475 3980 -425 3995
rect -475 3960 -460 3980
rect -440 3960 -425 3980
rect -475 3895 -425 3960
rect 85 3980 135 3995
rect 85 3960 100 3980
rect 120 3960 135 3980
rect -295 3910 -45 3925
rect -295 3895 -245 3910
rect -95 3895 -45 3910
rect 85 3895 135 3960
rect 185 3895 235 4025
rect 335 3935 385 3950
rect 335 3925 350 3935
rect 285 3915 350 3925
rect 370 3915 385 3935
rect 285 3905 385 3915
rect 285 3895 335 3905
rect -675 2680 -625 2695
rect -575 2680 -525 2695
rect -475 2680 -425 2695
rect -295 2655 -245 2695
rect -95 2655 -45 2695
rect 85 2680 135 2695
rect 185 2680 235 2695
rect 285 2680 335 2695
rect -730 2640 -45 2655
rect -625 2600 -575 2615
rect -525 2600 -475 2615
rect -425 2600 -375 2615
rect -325 2600 -275 2615
rect -65 2600 -15 2615
rect 35 2600 85 2615
rect 135 2600 185 2615
rect 235 2600 285 2615
rect -725 1370 -680 1385
rect -725 1350 -715 1370
rect -695 1355 -680 1370
rect -625 1375 -575 1400
rect -625 1355 -610 1375
rect -590 1355 -575 1375
rect -525 1385 -475 1400
rect -425 1385 -375 1400
rect -525 1355 -375 1385
rect -695 1350 -575 1355
rect -725 1340 -575 1350
rect -425 1315 -375 1355
rect -325 1385 -275 1400
rect -65 1385 -15 1400
rect -325 1375 -15 1385
rect -325 1355 -310 1375
rect -290 1355 -50 1375
rect -30 1355 -15 1375
rect -325 1340 -15 1355
rect 35 1385 85 1400
rect 135 1385 185 1400
rect 35 1355 185 1385
rect 235 1375 285 1400
rect 235 1355 250 1375
rect 270 1355 285 1375
rect 35 1315 85 1355
rect 235 1340 285 1355
rect -725 1305 85 1315
rect -725 1285 -715 1305
rect -695 1300 85 1305
rect -695 1285 -680 1300
rect -725 1270 -680 1285
rect -425 1260 -375 1275
rect -425 1240 -410 1260
rect -390 1240 -375 1260
rect -625 1215 -575 1230
rect -525 1215 -475 1230
rect -425 1215 -375 1240
rect 35 1260 85 1275
rect 35 1240 50 1260
rect 70 1240 85 1260
rect -325 1215 -275 1230
rect -65 1215 -15 1230
rect 35 1215 85 1240
rect 135 1215 185 1230
rect 235 1215 285 1230
rect -625 -20 -575 15
rect -525 5 -475 15
rect -425 5 -375 15
rect -525 -10 -375 5
rect -625 -40 -610 -20
rect -590 -40 -575 -20
rect -730 -55 -575 -40
rect -325 -20 -275 15
rect -325 -40 -310 -20
rect -290 -40 -275 -20
rect -325 -55 -275 -40
rect -65 -20 -15 15
rect 35 5 85 15
rect 135 5 185 15
rect 35 -10 185 5
rect -65 -40 -50 -20
rect -30 -40 -15 -20
rect -65 -55 -15 -40
rect 235 -20 285 15
rect 235 -40 250 -20
rect 270 -40 285 -20
rect 235 -55 285 -40
<< polycont >>
rect -710 3920 -690 3940
rect -460 3960 -440 3980
rect 100 3960 120 3980
rect 350 3915 370 3935
rect -715 1350 -695 1370
rect -610 1355 -590 1375
rect -310 1355 -290 1375
rect -50 1355 -30 1375
rect 250 1355 270 1375
rect -715 1285 -695 1305
rect -410 1240 -390 1260
rect 50 1240 70 1260
rect -610 -40 -590 -20
rect -310 -40 -290 -20
rect -50 -40 -30 -20
rect 250 -40 270 -20
<< locali >>
rect 85 3990 390 3995
rect -475 3980 390 3990
rect -475 3960 -460 3980
rect -440 3960 100 3980
rect 120 3970 390 3980
rect 120 3960 135 3970
rect -475 3950 135 3960
rect -725 3940 -675 3950
rect -725 3920 -710 3940
rect -690 3920 -675 3940
rect 335 3935 385 3945
rect -725 3910 -675 3920
rect -520 3910 180 3930
rect -720 3880 -680 3910
rect -720 2710 -710 3880
rect -690 2710 -680 3880
rect -720 2700 -680 2710
rect -620 3880 -580 3890
rect -620 2710 -610 3880
rect -590 2710 -580 3880
rect -620 2650 -580 2710
rect -520 3880 -480 3910
rect -520 2710 -510 3880
rect -490 2710 -480 3880
rect -520 2700 -480 2710
rect -420 3880 -380 3890
rect -420 2710 -410 3880
rect -390 2710 -380 3880
rect -420 2650 -380 2710
rect -340 3880 -300 3910
rect -340 2710 -330 3880
rect -310 2710 -300 3880
rect -340 2700 -300 2710
rect -240 3880 -100 3890
rect -240 2710 -230 3880
rect -210 2710 -180 3880
rect -160 2710 -130 3880
rect -110 2710 -100 3880
rect -240 2700 -100 2710
rect -40 3880 0 3910
rect -40 2710 -30 3880
rect -10 2710 0 3880
rect -40 2700 0 2710
rect 40 3880 80 3890
rect 40 2710 50 3880
rect 70 2710 80 3880
rect 40 2650 80 2710
rect 140 3880 180 3910
rect 335 3915 350 3935
rect 370 3915 385 3935
rect 335 3905 385 3915
rect 140 2710 150 3880
rect 170 2710 180 3880
rect 140 2700 180 2710
rect 240 3880 280 3890
rect 240 2710 250 3880
rect 270 2710 280 3880
rect 240 2650 280 2710
rect 340 3880 380 3905
rect 340 2710 350 3880
rect 370 2710 380 3880
rect 340 2700 380 2710
rect -620 2630 -530 2650
rect -670 2585 -630 2595
rect -670 1415 -660 2585
rect -640 1415 -630 2585
rect -670 1405 -630 1415
rect -570 2585 -530 2630
rect -420 2625 -330 2650
rect -570 1415 -560 2585
rect -540 1415 -530 2585
rect -570 1405 -530 1415
rect -470 2585 -430 2595
rect -470 1415 -460 2585
rect -440 1415 -430 2585
rect -470 1405 -430 1415
rect -370 2585 -330 2625
rect -10 2625 80 2650
rect 190 2625 280 2650
rect -370 1415 -360 2585
rect -340 1415 -330 2585
rect -370 1405 -330 1415
rect -270 2585 -230 2595
rect -270 1415 -260 2585
rect -240 1415 -230 2585
rect -270 1405 -230 1415
rect -190 2585 -150 2595
rect -190 1415 -180 2585
rect -160 1415 -150 2585
rect -190 1405 -150 1415
rect -110 2585 -70 2595
rect -110 1415 -100 2585
rect -80 1415 -70 2585
rect -110 1405 -70 1415
rect -10 2585 30 2625
rect -10 1415 0 2585
rect 20 1415 30 2585
rect -10 1405 30 1415
rect 90 2585 130 2595
rect 90 1415 100 2585
rect 120 1415 130 2585
rect 90 1405 130 1415
rect 190 2585 230 2625
rect 190 1415 200 2585
rect 220 1415 230 2585
rect 190 1405 230 1415
rect 290 2585 330 2595
rect 290 1415 300 2585
rect 320 1415 330 2585
rect 290 1405 330 1415
rect -725 1370 -680 1385
rect -725 1360 -715 1370
rect -730 1350 -715 1360
rect -695 1350 -680 1370
rect -730 1340 -680 1350
rect -725 1305 -680 1315
rect -725 1290 -715 1305
rect -730 1285 -715 1290
rect -695 1285 -680 1305
rect -730 1270 -680 1285
rect -660 1300 -640 1405
rect -620 1375 -280 1385
rect -620 1355 -610 1375
rect -590 1355 -310 1375
rect -290 1355 -280 1375
rect -620 1345 -280 1355
rect -660 1285 -560 1300
rect -660 1265 -645 1285
rect -575 1265 -560 1285
rect -260 1270 -230 1405
rect -110 1270 -80 1405
rect -60 1375 280 1385
rect -60 1355 -50 1375
rect -30 1355 250 1375
rect 270 1355 280 1375
rect -60 1345 280 1355
rect 300 1300 320 1405
rect 215 1290 320 1300
rect 215 1285 390 1290
rect -660 1250 -560 1265
rect -425 1260 85 1270
rect -660 1215 -640 1250
rect -425 1240 -410 1260
rect -390 1240 50 1260
rect 70 1240 85 1260
rect 215 1265 230 1285
rect 305 1265 390 1285
rect 215 1260 390 1265
rect 215 1250 320 1260
rect -425 1230 85 1240
rect -670 1210 -640 1215
rect -670 1200 -630 1210
rect -670 30 -660 1200
rect -640 30 -630 1200
rect -670 20 -630 30
rect -470 1200 -430 1210
rect -260 1205 -230 1230
rect -110 1210 -80 1230
rect 300 1210 320 1250
rect -470 30 -460 1200
rect -440 30 -430 1200
rect -470 20 -430 30
rect -270 1200 -230 1205
rect -270 30 -260 1200
rect -240 30 -230 1200
rect -270 20 -230 30
rect -195 1200 -150 1210
rect -195 30 -180 1200
rect -160 30 -150 1200
rect -195 20 -150 30
rect -110 1200 -70 1210
rect -110 30 -100 1200
rect -80 30 -70 1200
rect -110 20 -70 30
rect 90 1200 130 1210
rect 90 30 100 1200
rect 120 30 130 1200
rect 90 20 130 30
rect 290 1200 330 1210
rect 290 30 300 1200
rect 320 30 330 1200
rect 290 20 330 30
rect -625 -20 -575 -10
rect -625 -40 -610 -20
rect -590 -40 -575 -20
rect -625 -50 -575 -40
rect -325 -20 -275 -10
rect -325 -40 -310 -20
rect -290 -40 -275 -20
rect -325 -50 -275 -40
rect -65 -20 -15 -10
rect -65 -40 -50 -20
rect -30 -40 -15 -20
rect -65 -50 -15 -40
rect 235 -20 285 -10
rect 235 -40 250 -20
rect 270 -40 285 -20
rect 235 -50 285 -40
<< viali >>
rect -710 2710 -690 3880
rect -230 2710 -210 3880
rect -180 2710 -160 3880
rect -130 2710 -110 3880
rect 350 2710 370 3880
rect -460 1415 -440 2585
rect -180 1415 -160 2585
rect 100 1415 120 2585
rect -645 1265 -575 1285
rect 230 1265 305 1285
rect -460 30 -440 1200
rect -180 30 -160 1200
rect 100 30 120 1200
rect -610 -40 -590 -20
rect -310 -40 -290 -20
rect -50 -40 -30 -20
rect 250 -40 270 -20
<< metal1 >>
rect -730 3880 390 3890
rect -730 2710 -710 3880
rect -690 2710 -230 3880
rect -210 2710 -180 3880
rect -160 2710 -130 3880
rect -110 2710 350 3880
rect 370 2710 390 3880
rect -730 2700 390 2710
rect -225 2595 -195 2600
rect -730 2585 390 2595
rect -730 1415 -460 2585
rect -440 1415 -180 2585
rect -160 1415 100 2585
rect 120 1415 390 2585
rect -730 1405 390 1415
rect -225 1400 -195 1405
rect -660 1285 320 1300
rect -660 1265 -645 1285
rect -575 1265 230 1285
rect 305 1265 320 1285
rect -660 1250 320 1265
rect -730 1200 390 1210
rect -730 30 -460 1200
rect -440 30 -180 1200
rect -160 30 100 1200
rect 120 30 390 1200
rect -730 20 390 30
rect -625 -20 285 -10
rect -625 -40 -610 -20
rect -590 -40 -310 -20
rect -290 -40 -50 -20
rect -30 -40 250 -20
rect 270 -40 285 -20
rect -625 -55 285 -40
<< labels >>
rlabel metal1 -730 2000 -730 2000 7 VP
port 9 w
rlabel poly -730 -45 -730 -45 7 Vcn
port 6 w
rlabel metal1 -730 610 -730 610 7 VN
port 10 w
rlabel poly -730 2645 -730 2645 7 Vbn
port 1 w
rlabel metal1 -730 3295 -730 3295 7 VN
port 8 w
rlabel poly 390 4030 390 4030 3 Vref
port 3 w
rlabel locali -730 1350 -730 1350 7 Vcp
port 5 w
rlabel locali 390 1275 390 1275 3 Vout
port 7 e
rlabel locali 390 3985 390 3985 3 Vin
port 2 e
rlabel locali -730 1280 -730 1280 7 Vbp
port 4 w
<< end >>
