magic
tech sky130A
timestamp 1698126361
<< nwell >>
rect -830 1360 490 2610
<< nmos >>
rect -775 2695 -725 3895
rect -675 2695 -625 3895
rect -575 2695 -525 3895
rect -475 2695 -425 3895
rect -295 2695 -245 3895
rect -95 2695 -45 3895
rect 85 2695 135 3895
rect 185 2695 235 3895
rect 285 2695 335 3895
rect 385 2695 435 3895
rect -725 0 -675 1200
rect -625 0 -575 1200
rect -525 0 -475 1200
rect -425 0 -375 1200
rect -325 0 -275 1200
rect -65 0 -15 1200
rect 35 0 85 1200
rect 135 0 185 1200
rect 235 0 285 1200
rect 335 0 385 1200
<< pmos >>
rect -725 1385 -675 2585
rect -625 1385 -575 2585
rect -525 1385 -475 2585
rect -425 1385 -375 2585
rect -325 1385 -275 2585
rect -65 1385 -15 2585
rect 35 1385 85 2585
rect 135 1385 185 2585
rect 235 1385 285 2585
rect 335 1385 385 2585
<< ndiff >>
rect -825 3880 -775 3895
rect -825 2710 -810 3880
rect -790 2710 -775 3880
rect -825 2695 -775 2710
rect -725 3880 -675 3895
rect -725 2710 -710 3880
rect -690 2710 -675 3880
rect -725 2695 -675 2710
rect -625 3880 -575 3895
rect -625 2710 -610 3880
rect -590 2710 -575 3880
rect -625 2695 -575 2710
rect -525 3880 -475 3895
rect -525 2710 -510 3880
rect -490 2710 -475 3880
rect -525 2695 -475 2710
rect -425 3880 -375 3895
rect -425 2710 -410 3880
rect -390 2710 -375 3880
rect -425 2695 -375 2710
rect -345 3880 -295 3895
rect -345 2710 -330 3880
rect -310 2710 -295 3880
rect -345 2695 -295 2710
rect -245 3880 -195 3895
rect -145 3880 -95 3895
rect -245 2710 -230 3880
rect -210 2710 -195 3880
rect -145 2710 -130 3880
rect -110 2710 -95 3880
rect -245 2695 -195 2710
rect -145 2695 -95 2710
rect -45 3880 5 3895
rect -45 2710 -30 3880
rect -10 2710 5 3880
rect -45 2695 5 2710
rect 35 3880 85 3895
rect 35 2710 50 3880
rect 70 2710 85 3880
rect 35 2695 85 2710
rect 135 3880 185 3895
rect 135 2710 150 3880
rect 170 2710 185 3880
rect 135 2695 185 2710
rect 235 3880 285 3895
rect 235 2710 250 3880
rect 270 2710 285 3880
rect 235 2695 285 2710
rect 335 3880 385 3895
rect 335 2710 350 3880
rect 370 2710 385 3880
rect 335 2695 385 2710
rect 435 3880 485 3895
rect 435 2710 450 3880
rect 470 2710 485 3880
rect 435 2695 485 2710
rect -775 1185 -725 1200
rect -775 15 -760 1185
rect -740 15 -725 1185
rect -775 0 -725 15
rect -675 1185 -625 1200
rect -675 15 -660 1185
rect -640 15 -625 1185
rect -675 0 -625 15
rect -575 0 -525 1200
rect -475 1185 -425 1200
rect -475 15 -460 1185
rect -440 15 -425 1185
rect -475 0 -425 15
rect -375 0 -325 1200
rect -275 1185 -225 1200
rect -275 15 -260 1185
rect -240 15 -225 1185
rect -275 0 -225 15
rect -115 1185 -65 1200
rect -115 15 -100 1185
rect -80 15 -65 1185
rect -115 0 -65 15
rect -15 0 35 1200
rect 85 1185 135 1200
rect 85 15 100 1185
rect 120 15 135 1185
rect 85 0 135 15
rect 185 0 235 1200
rect 285 1185 335 1200
rect 285 15 300 1185
rect 320 15 335 1185
rect 285 0 335 15
rect 385 1185 435 1200
rect 385 15 400 1185
rect 420 15 435 1185
rect 385 0 435 15
<< pdiff >>
rect -775 2570 -725 2585
rect -775 1400 -760 2570
rect -740 1400 -725 2570
rect -775 1385 -725 1400
rect -675 2570 -625 2585
rect -675 1400 -660 2570
rect -640 1400 -625 2570
rect -675 1385 -625 1400
rect -575 2570 -525 2585
rect -575 1400 -560 2570
rect -540 1400 -525 2570
rect -575 1385 -525 1400
rect -475 2570 -425 2585
rect -475 1400 -460 2570
rect -440 1400 -425 2570
rect -475 1385 -425 1400
rect -375 2570 -325 2585
rect -375 1400 -360 2570
rect -340 1400 -325 2570
rect -375 1385 -325 1400
rect -275 2570 -225 2585
rect -275 1400 -260 2570
rect -240 1400 -225 2570
rect -275 1390 -225 1400
rect -275 1385 -230 1390
rect -115 2570 -65 2585
rect -115 1400 -100 2570
rect -80 1400 -65 2570
rect -115 1385 -65 1400
rect -15 2570 35 2585
rect -15 1400 0 2570
rect 20 1400 35 2570
rect -15 1385 35 1400
rect 85 2570 135 2585
rect 85 1400 100 2570
rect 120 1400 135 2570
rect 85 1385 135 1400
rect 185 2570 235 2585
rect 185 1400 200 2570
rect 220 1400 235 2570
rect 185 1385 235 1400
rect 285 2570 335 2585
rect 285 1400 300 2570
rect 320 1400 335 2570
rect 285 1385 335 1400
rect 385 2570 435 2585
rect 385 1400 400 2570
rect 420 1400 435 2570
rect 385 1385 435 1400
<< ndiffc >>
rect -810 2710 -790 3880
rect -710 2710 -690 3880
rect -610 2710 -590 3880
rect -510 2710 -490 3880
rect -410 2710 -390 3880
rect -330 2710 -310 3880
rect -230 2710 -210 3880
rect -130 2710 -110 3880
rect -30 2710 -10 3880
rect 50 2710 70 3880
rect 150 2710 170 3880
rect 250 2710 270 3880
rect 350 2710 370 3880
rect 450 2710 470 3880
rect -760 15 -740 1185
rect -660 15 -640 1185
rect -460 15 -440 1185
rect -260 15 -240 1185
rect -100 15 -80 1185
rect 100 15 120 1185
rect 300 15 320 1185
rect 400 15 420 1185
<< pdiffc >>
rect -760 1400 -740 2570
rect -660 1400 -640 2570
rect -560 1400 -540 2570
rect -460 1400 -440 2570
rect -360 1400 -340 2570
rect -260 1400 -240 2570
rect -100 1400 -80 2570
rect 0 1400 20 2570
rect 100 1400 120 2570
rect 200 1400 220 2570
rect 300 1400 320 2570
rect 400 1400 420 2570
<< psubdiff >>
rect -195 3880 -145 3895
rect -195 2710 -180 3880
rect -160 2710 -145 3880
rect -195 2695 -145 2710
rect -195 1185 -145 1200
rect -195 15 -180 1185
rect -160 15 -145 1185
rect -195 0 -145 15
<< nsubdiff >>
rect -195 2570 -145 2585
rect -195 1400 -180 2570
rect -160 1400 -145 2570
rect -195 1385 -145 1400
<< psubdiffcont >>
rect -180 2710 -160 3880
rect -180 15 -160 1185
<< nsubdiffcont >>
rect -180 1400 -160 2570
<< poly >>
rect -575 4025 490 4040
rect -725 3940 -675 3955
rect -725 3925 -710 3940
rect -775 3920 -710 3925
rect -690 3925 -675 3940
rect -690 3920 -625 3925
rect -775 3910 -625 3920
rect -775 3895 -725 3910
rect -675 3895 -625 3910
rect -575 3895 -525 4025
rect -475 3980 -425 3995
rect -475 3960 -460 3980
rect -440 3960 -425 3980
rect -475 3895 -425 3960
rect 85 3980 135 3995
rect 85 3960 100 3980
rect 120 3960 135 3980
rect -295 3895 -245 3910
rect -95 3895 -45 3910
rect 85 3895 135 3960
rect 185 3895 235 4025
rect 335 3935 385 3950
rect 335 3925 350 3935
rect 285 3915 350 3925
rect 370 3925 385 3935
rect 370 3915 435 3925
rect 285 3905 435 3915
rect 285 3895 335 3905
rect 385 3895 435 3905
rect -775 2680 -725 2695
rect -675 2680 -625 2695
rect -575 2680 -525 2695
rect -475 2680 -425 2695
rect -295 2655 -245 2695
rect -95 2655 -45 2695
rect 85 2680 135 2695
rect 185 2680 235 2695
rect 285 2680 335 2695
rect 385 2680 435 2695
rect -830 2640 -45 2655
rect 385 2630 435 2645
rect 385 2620 400 2630
rect -830 2600 -675 2615
rect 335 2610 400 2620
rect 420 2610 435 2630
rect -830 2580 -820 2600
rect -800 2580 -785 2600
rect -725 2585 -675 2600
rect -625 2585 -575 2600
rect -525 2585 -475 2600
rect -425 2585 -375 2600
rect -325 2585 -275 2600
rect -65 2585 -15 2600
rect 35 2585 85 2600
rect 135 2585 185 2600
rect 235 2585 285 2600
rect 335 2595 435 2610
rect 335 2585 385 2595
rect -830 2565 -785 2580
rect -725 1370 -675 1385
rect -800 1355 -750 1370
rect -800 1335 -785 1355
rect -765 1340 -750 1355
rect -625 1360 -575 1385
rect -625 1340 -610 1360
rect -590 1340 -575 1360
rect -525 1370 -475 1385
rect -425 1370 -375 1385
rect -525 1340 -375 1370
rect -765 1335 -575 1340
rect -800 1325 -575 1335
rect -800 1320 -750 1325
rect -425 1300 -375 1340
rect -325 1370 -275 1385
rect -65 1370 -15 1385
rect -325 1360 -15 1370
rect -325 1340 -310 1360
rect -290 1340 -50 1360
rect -30 1340 -15 1360
rect -325 1325 -15 1340
rect 35 1370 85 1385
rect 135 1370 185 1385
rect 35 1340 185 1370
rect 235 1360 285 1385
rect 335 1370 385 1385
rect 235 1340 250 1360
rect 270 1340 285 1360
rect 35 1300 85 1340
rect 235 1325 285 1340
rect -730 1285 85 1300
rect -730 1265 -715 1285
rect -695 1265 -680 1285
rect -825 1245 -775 1260
rect -730 1255 -680 1265
rect -825 1225 -810 1245
rect -790 1225 -775 1245
rect -425 1245 -375 1260
rect -425 1225 -410 1245
rect -390 1225 -375 1245
rect -825 1210 -675 1225
rect -725 1200 -675 1210
rect -625 1200 -575 1215
rect -525 1200 -475 1215
rect -425 1200 -375 1225
rect 35 1245 85 1260
rect 35 1225 50 1245
rect 70 1225 85 1245
rect 385 1245 435 1260
rect 385 1230 400 1245
rect -325 1200 -275 1215
rect -65 1200 -15 1215
rect 35 1200 85 1225
rect 335 1225 400 1230
rect 420 1225 435 1245
rect 335 1215 435 1225
rect 135 1200 185 1215
rect 235 1200 285 1215
rect 335 1200 385 1215
rect -725 -15 -675 0
rect -625 -35 -575 0
rect -525 -10 -475 0
rect -425 -10 -375 0
rect -525 -25 -375 -10
rect -625 -55 -610 -35
rect -590 -55 -575 -35
rect -830 -70 -575 -55
rect -325 -35 -275 0
rect -325 -55 -310 -35
rect -290 -55 -275 -35
rect -325 -70 -275 -55
rect -65 -35 -15 0
rect 35 -10 85 0
rect 135 -10 185 0
rect 35 -25 185 -10
rect -65 -55 -50 -35
rect -30 -55 -15 -35
rect -65 -70 -15 -55
rect 235 -35 285 0
rect 335 -15 385 0
rect 235 -55 250 -35
rect 270 -55 285 -35
rect 235 -70 285 -55
<< polycont >>
rect -710 3920 -690 3940
rect -460 3960 -440 3980
rect 100 3960 120 3980
rect 350 3915 370 3935
rect 400 2610 420 2630
rect -820 2580 -800 2600
rect -785 1335 -765 1355
rect -610 1340 -590 1360
rect -310 1340 -290 1360
rect -50 1340 -30 1360
rect 250 1340 270 1360
rect -715 1265 -695 1285
rect -810 1225 -790 1245
rect -410 1225 -390 1245
rect 50 1225 70 1245
rect 400 1225 420 1245
rect -610 -55 -590 -35
rect -310 -55 -290 -35
rect -50 -55 -30 -35
rect 250 -55 270 -35
<< locali >>
rect 85 3990 490 3995
rect -475 3980 490 3990
rect -475 3960 -460 3980
rect -440 3960 100 3980
rect 120 3970 490 3980
rect 120 3960 135 3970
rect -475 3950 135 3960
rect -725 3940 -675 3950
rect -725 3920 -710 3940
rect -690 3920 -675 3940
rect 335 3935 385 3945
rect -725 3910 -675 3920
rect -520 3910 -300 3930
rect -820 3880 -780 3890
rect -820 2710 -810 3880
rect -790 2710 -780 3880
rect -820 2680 -780 2710
rect -720 3880 -680 3910
rect -720 2710 -710 3880
rect -690 2710 -680 3880
rect -720 2700 -680 2710
rect -620 3880 -580 3890
rect -620 2710 -610 3880
rect -590 2710 -580 3880
rect -820 2655 -645 2680
rect -830 2600 -730 2615
rect -830 2580 -820 2600
rect -800 2580 -730 2600
rect -830 2570 -730 2580
rect -830 2565 -760 2570
rect -770 1400 -760 2565
rect -740 1400 -730 2570
rect -770 1390 -730 1400
rect -670 2580 -645 2655
rect -620 2650 -580 2710
rect -520 3880 -480 3910
rect -520 2710 -510 3880
rect -490 2710 -480 3880
rect -520 2700 -480 2710
rect -420 3880 -380 3890
rect -420 2710 -410 3880
rect -390 2710 -380 3880
rect -420 2650 -380 2710
rect -340 3880 -300 3910
rect -40 3910 180 3930
rect -340 2710 -330 3880
rect -310 2710 -300 3880
rect -340 2700 -300 2710
rect -240 3880 -100 3890
rect -240 2710 -230 3880
rect -210 2710 -180 3880
rect -160 2710 -130 3880
rect -110 2710 -100 3880
rect -240 2700 -100 2710
rect -40 3880 0 3910
rect -40 2710 -30 3880
rect -10 2710 0 3880
rect -40 2700 0 2710
rect 40 3880 80 3890
rect 40 2710 50 3880
rect 70 2710 80 3880
rect 40 2650 80 2710
rect 140 3880 180 3910
rect 335 3915 350 3935
rect 370 3915 385 3935
rect 335 3905 385 3915
rect 140 2710 150 3880
rect 170 2710 180 3880
rect 140 2700 180 2710
rect 240 3880 280 3890
rect 240 2710 250 3880
rect 270 2710 280 3880
rect 240 2650 280 2710
rect 340 3880 380 3905
rect 340 2710 350 3880
rect 370 2710 380 3880
rect 340 2700 380 2710
rect 440 3880 480 3890
rect 440 2710 450 3880
rect 470 2710 480 3880
rect 440 2680 480 2710
rect -620 2625 -530 2650
rect -420 2625 -330 2650
rect -670 2570 -630 2580
rect -670 1400 -660 2570
rect -640 1400 -630 2570
rect -670 1390 -630 1400
rect -570 2570 -530 2625
rect -570 1400 -560 2570
rect -540 1400 -530 2570
rect -570 1390 -530 1400
rect -470 2570 -430 2580
rect -470 1400 -460 2570
rect -440 1400 -430 2570
rect -470 1390 -430 1400
rect -370 2570 -330 2625
rect -10 2625 80 2650
rect 190 2625 280 2650
rect 305 2660 480 2680
rect -370 1400 -360 2570
rect -340 1400 -330 2570
rect -370 1390 -330 1400
rect -270 2570 -230 2580
rect -270 1400 -260 2570
rect -240 1400 -230 2570
rect -270 1390 -230 1400
rect -190 2570 -150 2580
rect -190 1400 -180 2570
rect -160 1400 -150 2570
rect -190 1390 -150 1400
rect -110 2570 -70 2580
rect -110 1400 -100 2570
rect -80 1400 -70 2570
rect -110 1390 -70 1400
rect -10 2570 30 2625
rect -10 1400 0 2570
rect 20 1400 30 2570
rect -10 1390 30 1400
rect 90 2570 130 2580
rect 90 1400 100 2570
rect 120 1400 130 2570
rect 90 1390 130 1400
rect 190 2570 230 2625
rect 305 2580 330 2660
rect 385 2630 435 2640
rect 385 2610 400 2630
rect 420 2610 435 2630
rect 385 2595 435 2610
rect 190 1400 200 2570
rect 220 1400 230 2570
rect 190 1390 230 1400
rect 290 2570 330 2580
rect 290 1400 300 2570
rect 320 1400 330 2570
rect 290 1390 330 1400
rect 390 2570 430 2595
rect 390 1400 400 2570
rect 420 1400 430 2570
rect 390 1390 430 1400
rect -800 1355 -750 1370
rect -800 1345 -785 1355
rect -830 1335 -785 1345
rect -765 1335 -750 1355
rect -830 1325 -750 1335
rect -800 1320 -750 1325
rect -830 1285 -680 1300
rect -830 1280 -715 1285
rect -730 1265 -715 1280
rect -695 1265 -680 1285
rect -825 1245 -775 1260
rect -730 1255 -680 1265
rect -825 1225 -810 1245
rect -790 1235 -775 1245
rect -790 1225 -730 1235
rect -825 1210 -730 1225
rect -770 1185 -730 1210
rect -660 1195 -640 1390
rect -620 1360 -280 1370
rect -620 1340 -610 1360
rect -590 1340 -310 1360
rect -290 1340 -280 1360
rect -620 1330 -280 1340
rect -260 1255 -230 1390
rect -110 1255 -80 1390
rect -60 1360 280 1370
rect -60 1340 -50 1360
rect -30 1340 250 1360
rect 270 1340 280 1360
rect -60 1330 280 1340
rect 300 1355 320 1390
rect 300 1325 490 1355
rect -425 1245 85 1255
rect -425 1225 -410 1245
rect -390 1225 50 1245
rect 70 1225 85 1245
rect -425 1215 85 1225
rect -260 1195 -230 1215
rect -110 1195 -80 1215
rect 300 1195 320 1325
rect 385 1245 435 1260
rect 385 1225 400 1245
rect 420 1225 435 1245
rect 385 1215 435 1225
rect -770 15 -760 1185
rect -740 15 -730 1185
rect -770 5 -730 15
rect -670 1185 -630 1195
rect -670 15 -660 1185
rect -640 15 -630 1185
rect -670 5 -630 15
rect -470 1185 -430 1195
rect -470 15 -460 1185
rect -440 15 -430 1185
rect -470 5 -430 15
rect -270 1185 -230 1195
rect -270 15 -260 1185
rect -240 15 -230 1185
rect -270 5 -230 15
rect -190 1185 -150 1195
rect -190 15 -180 1185
rect -160 15 -150 1185
rect -190 5 -150 15
rect -110 1185 -70 1195
rect -110 15 -100 1185
rect -80 15 -70 1185
rect -110 5 -70 15
rect 90 1185 130 1195
rect 90 15 100 1185
rect 120 15 130 1185
rect 90 5 130 15
rect 290 1185 330 1195
rect 290 15 300 1185
rect 320 15 330 1185
rect 290 5 330 15
rect 390 1185 430 1215
rect 390 15 400 1185
rect 420 15 430 1185
rect 390 5 430 15
rect -625 -35 -575 -25
rect -625 -55 -610 -35
rect -590 -55 -575 -35
rect -625 -65 -575 -55
rect -325 -35 -275 -25
rect -325 -55 -310 -35
rect -290 -55 -275 -35
rect -325 -65 -275 -55
rect -65 -35 -15 -25
rect -65 -55 -50 -35
rect -30 -55 -15 -35
rect -65 -65 -15 -55
rect 235 -35 285 -25
rect 235 -55 250 -35
rect 270 -55 285 -35
rect 235 -65 285 -55
<< viali >>
rect -710 2710 -690 3880
rect -760 1400 -740 2570
rect -230 2710 -210 3880
rect -180 2710 -160 3880
rect -130 2710 -110 3880
rect 350 2710 370 3880
rect -460 1400 -440 2570
rect -180 1400 -160 2570
rect 100 1400 120 2570
rect 400 1400 420 2570
rect -760 15 -740 1185
rect -460 15 -440 1185
rect -180 15 -160 1185
rect 100 15 120 1185
rect 400 15 420 1185
rect -610 -55 -590 -35
rect -310 -55 -290 -35
rect -50 -55 -30 -35
rect 250 -55 270 -35
<< metal1 >>
rect 385 3890 435 3895
rect -830 3880 490 3890
rect -830 2710 -710 3880
rect -690 2710 -230 3880
rect -210 2710 -180 3880
rect -160 2710 -130 3880
rect -110 2710 350 3880
rect 370 2710 490 3880
rect -830 2700 490 2710
rect 385 2695 435 2700
rect -830 2570 490 2580
rect -830 1400 -760 2570
rect -740 1400 -460 2570
rect -440 1400 -180 2570
rect -160 1400 100 2570
rect 120 1400 400 2570
rect 420 1400 490 2570
rect -830 1390 490 1400
rect -830 1185 490 1195
rect -830 15 -760 1185
rect -740 15 -460 1185
rect -440 15 -180 1185
rect -160 15 100 1185
rect 120 15 400 1185
rect 420 15 490 1185
rect -830 5 490 15
rect -625 -35 285 -25
rect -625 -55 -610 -35
rect -590 -55 -310 -35
rect -290 -55 -50 -35
rect -30 -55 250 -35
rect 270 -55 285 -35
rect -625 -70 285 -55
<< labels >>
rlabel poly -830 2645 -830 2645 7 Vbn
port 1 w
rlabel metal1 -830 3295 -830 3295 7 VN
port 8 w
rlabel poly 490 4030 490 4030 3 Vref
port 3 w
rlabel locali 490 3985 490 3985 3 Vin
port 2 e
rlabel locali 490 1340 490 1340 3 Vout
port 7 e
rlabel locali -830 1290 -830 1290 7 Vbp
port 4 w
rlabel metal1 -830 1985 -830 1985 7 VP
port 9 w
rlabel poly -830 -60 -830 -60 7 Vcn
port 6 w
rlabel metal1 -830 595 -830 595 7 VN
port 10 w
rlabel locali -830 1335 -830 1335 7 Vcp
port 5 w
<< end >>
