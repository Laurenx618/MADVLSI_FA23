magic
tech sky130A
timestamp 1698134376
<< poly >>
rect 3240 4390 3290 4405
rect 1930 3005 2030 3020
rect 1930 2610 1945 3005
rect 1940 310 1955 1285
rect 1940 295 2060 310
<< locali >>
rect 3240 4335 3290 4360
rect 1940 1710 1960 2620
rect 1940 1690 2015 1710
rect 3240 1690 3290 1720
rect 1935 1645 2015 1665
rect 1935 1255 1955 1645
<< metal1 >>
rect -10 3975 10 5165
rect 1920 3975 1940 5165
rect -10 1365 10 3865
rect 1970 3065 1990 4255
rect 3270 3065 3290 4255
rect 1970 2715 1990 2945
rect 1970 1755 1990 2605
rect 3270 1755 3290 2945
rect -10 65 10 1255
rect 1920 65 1940 1255
rect 1970 370 1990 1560
rect 3270 370 3290 1560
use diff_amp  diff_amp_0
timestamp 1698126361
transform 1 0 2800 0 1 365
box -830 -70 490 4040
use v_gen  v_gen_0
timestamp 1698134288
transform 1 0 360 0 1 2530
box -370 -2560 1580 2675
<< labels >>
rlabel metal1 -10 4580 -10 4580 7 VP
rlabel metal1 -10 660 -10 660 7 VP
rlabel metal1 1970 2350 1970 2350 7 VP
rlabel metal1 -10 2610 -10 2610 7 VN
rlabel metal1 1970 960 1970 960 7 VN
rlabel metal1 1970 3660 1970 3660 7 VN
rlabel poly 3290 4395 3290 4395 3 Vref
rlabel locali 3290 4350 3290 4350 3 Vin
rlabel locali 3290 1705 3290 1705 3 Vout
<< end >>
