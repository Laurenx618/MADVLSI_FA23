magic
tech sky130A
timestamp 1694896595
<< nwell >>
rect -100 345 455 705
<< nmos >>
rect -20 150 -5 250
rect 20 150 35 250
rect 85 150 100 250
rect 235 150 250 250
rect 300 150 315 250
rect 365 150 380 250
rect -20 -65 -5 35
rect 20 -65 35 35
rect 85 -65 100 35
rect 235 -65 250 35
rect 300 -65 315 35
rect 365 -65 380 35
<< pmos >>
rect -20 585 -5 685
rect 45 585 60 685
rect 110 585 125 685
rect 260 585 275 685
rect 300 585 315 685
rect 365 585 380 685
rect -20 370 -5 470
rect 45 370 60 470
rect 110 370 125 470
rect 260 370 275 470
rect 300 370 315 470
rect 365 370 380 470
<< ndiff >>
rect -70 235 -20 250
rect -70 165 -55 235
rect -35 165 -20 235
rect -70 150 -20 165
rect -5 150 20 250
rect 35 235 85 250
rect 35 165 50 235
rect 70 165 85 235
rect 35 150 85 165
rect 100 235 150 250
rect 100 165 115 235
rect 135 165 150 235
rect 100 150 150 165
rect 185 235 235 250
rect 185 165 200 235
rect 220 165 235 235
rect 185 150 235 165
rect 250 235 300 250
rect 250 165 265 235
rect 285 165 300 235
rect 250 150 300 165
rect 315 235 365 250
rect 315 165 330 235
rect 350 165 365 235
rect 315 150 365 165
rect 380 235 430 250
rect 380 165 395 235
rect 415 165 430 235
rect 380 150 430 165
rect -70 20 -20 35
rect -70 -50 -55 20
rect -35 -50 -20 20
rect -70 -65 -20 -50
rect -5 -65 20 35
rect 35 20 85 35
rect 35 -50 50 20
rect 70 -50 85 20
rect 35 -65 85 -50
rect 100 20 150 35
rect 100 -50 115 20
rect 135 -50 150 20
rect 100 -65 150 -50
rect 185 20 235 35
rect 185 -50 200 20
rect 220 -50 235 20
rect 185 -65 235 -50
rect 250 20 300 35
rect 250 -50 265 20
rect 285 -50 300 20
rect 250 -65 300 -50
rect 315 20 365 35
rect 315 -50 330 20
rect 350 -50 365 20
rect 315 -65 365 -50
rect 380 20 430 35
rect 380 -50 395 20
rect 415 -50 430 20
rect 380 -65 430 -50
<< pdiff >>
rect -70 670 -20 685
rect -70 600 -55 670
rect -35 600 -20 670
rect -70 585 -20 600
rect -5 670 45 685
rect -5 600 10 670
rect 30 600 45 670
rect -5 585 45 600
rect 60 670 110 685
rect 60 600 75 670
rect 95 600 110 670
rect 60 585 110 600
rect 125 670 175 685
rect 125 600 140 670
rect 160 600 175 670
rect 125 585 175 600
rect 210 670 260 685
rect 210 600 225 670
rect 245 600 260 670
rect 210 585 260 600
rect 275 585 300 685
rect 315 670 365 685
rect 315 600 330 670
rect 350 600 365 670
rect 315 585 365 600
rect 380 670 430 685
rect 380 600 395 670
rect 415 600 430 670
rect 380 585 430 600
rect -70 455 -20 470
rect -70 385 -55 455
rect -35 385 -20 455
rect -70 370 -20 385
rect -5 455 45 470
rect -5 385 10 455
rect 30 385 45 455
rect -5 370 45 385
rect 60 455 110 470
rect 60 385 75 455
rect 95 385 110 455
rect 60 370 110 385
rect 125 455 175 470
rect 125 385 140 455
rect 160 385 175 455
rect 125 370 175 385
rect 210 455 260 470
rect 210 385 225 455
rect 245 385 260 455
rect 210 370 260 385
rect 275 370 300 470
rect 315 455 365 470
rect 315 385 330 455
rect 350 385 365 455
rect 315 370 365 385
rect 380 455 430 470
rect 380 385 395 455
rect 415 385 430 455
rect 380 370 430 385
<< ndiffc >>
rect -55 165 -35 235
rect 50 165 70 235
rect 115 165 135 235
rect 200 165 220 235
rect 265 165 285 235
rect 330 165 350 235
rect 395 165 415 235
rect -55 -50 -35 20
rect 50 -50 70 20
rect 115 -50 135 20
rect 200 -50 220 20
rect 265 -50 285 20
rect 330 -50 350 20
rect 395 -50 415 20
<< pdiffc >>
rect -55 600 -35 670
rect 10 600 30 670
rect 75 600 95 670
rect 140 600 160 670
rect 225 600 245 670
rect 330 600 350 670
rect 395 600 415 670
rect -55 385 -35 455
rect 10 385 30 455
rect 75 385 95 455
rect 140 385 160 455
rect 225 385 245 455
rect 330 385 350 455
rect 395 385 415 455
<< psubdiff >>
rect 185 105 285 120
rect 185 85 200 105
rect 270 85 285 105
rect 185 70 285 85
<< nsubdiff >>
rect -70 535 30 550
rect -70 515 -55 535
rect 15 515 30 535
rect -70 500 30 515
<< psubdiffcont >>
rect 200 85 270 105
<< nsubdiffcont >>
rect -55 515 15 535
<< poly >>
rect 340 730 380 740
rect 340 710 350 730
rect 370 710 380 730
rect 340 700 380 710
rect -20 685 -5 700
rect 45 685 60 700
rect 110 685 125 700
rect 260 685 275 700
rect 300 685 315 700
rect 365 685 380 700
rect -20 575 -5 585
rect -80 560 -5 575
rect -20 470 -5 485
rect 45 470 60 585
rect 110 570 125 585
rect 260 570 275 585
rect 85 555 125 570
rect 85 535 95 555
rect 115 535 125 555
rect 85 525 125 535
rect 150 555 275 570
rect 150 535 160 555
rect 180 550 275 555
rect 180 535 190 550
rect 150 525 190 535
rect 150 500 165 525
rect 110 485 165 500
rect 110 470 125 485
rect 260 470 275 485
rect 300 470 315 585
rect 365 570 380 585
rect 405 560 455 575
rect 405 525 420 560
rect 340 515 420 525
rect 340 495 350 515
rect 370 510 420 515
rect 370 495 380 510
rect 340 485 380 495
rect 365 470 380 485
rect -20 310 -5 370
rect 45 360 60 370
rect 110 360 125 370
rect -45 300 -5 310
rect -45 280 -35 300
rect -15 280 -5 300
rect -45 270 -5 280
rect -20 250 -5 270
rect 20 345 60 360
rect 85 345 125 360
rect 260 355 275 370
rect 235 345 275 355
rect 20 250 35 345
rect 85 250 100 345
rect 235 325 245 345
rect 265 325 275 345
rect 235 315 275 325
rect 235 250 250 315
rect 300 250 315 370
rect 365 250 380 370
rect -20 135 -5 150
rect -80 45 -5 60
rect -20 35 -5 45
rect 20 35 35 150
rect 85 135 100 150
rect 235 135 250 150
rect 60 125 100 135
rect 60 105 70 125
rect 90 110 100 125
rect 90 105 140 110
rect 60 95 140 105
rect 125 60 140 95
rect 85 35 100 50
rect 125 45 250 60
rect 235 35 250 45
rect 300 35 315 150
rect 365 140 380 150
rect 365 125 420 140
rect 340 80 380 90
rect 340 60 350 80
rect 370 60 380 80
rect 340 50 380 60
rect 365 35 380 50
rect 405 85 420 125
rect 405 75 445 85
rect 405 55 415 75
rect 435 55 445 75
rect 405 45 445 55
rect -20 -80 -5 -65
rect 20 -120 35 -65
rect 85 -80 100 -65
rect 235 -80 250 -65
rect 300 -80 315 -65
rect 60 -90 100 -80
rect 60 -110 70 -90
rect 90 -110 100 -90
rect 60 -120 100 -110
rect 365 -120 380 -65
rect -5 -130 35 -120
rect -5 -150 5 -130
rect 25 -150 35 -130
rect -5 -160 35 -150
rect 340 -130 380 -120
rect 340 -150 350 -130
rect 370 -150 380 -130
rect 340 -160 380 -150
<< polycont >>
rect 350 710 370 730
rect 95 535 115 555
rect 160 535 180 555
rect 350 495 370 515
rect -35 280 -15 300
rect 245 325 265 345
rect 70 105 90 125
rect 350 60 370 80
rect 415 55 435 75
rect 70 -110 90 -90
rect 5 -150 25 -130
rect 350 -150 370 -130
<< locali >>
rect 340 730 380 740
rect -45 705 85 725
rect 340 720 350 730
rect -45 680 -25 705
rect 65 680 85 705
rect 280 710 350 720
rect 370 710 380 730
rect 280 700 380 710
rect -65 670 -25 680
rect -65 600 -55 670
rect -35 600 -25 670
rect -65 590 -25 600
rect 0 670 40 680
rect 0 600 10 670
rect 30 600 40 670
rect 0 590 40 600
rect 65 670 105 680
rect 65 600 75 670
rect 95 600 105 670
rect 65 590 105 600
rect 130 670 170 680
rect 130 600 140 670
rect 160 600 170 670
rect 130 590 170 600
rect 0 545 20 590
rect 150 570 170 590
rect 215 670 255 680
rect 215 600 225 670
rect 245 600 255 670
rect 215 590 255 600
rect 85 555 125 570
rect -65 535 25 545
rect -65 515 -55 535
rect 15 515 25 535
rect 85 535 95 555
rect 115 535 125 555
rect 85 525 125 535
rect 150 555 190 570
rect 150 535 160 555
rect 180 535 190 555
rect 150 525 190 535
rect -65 505 25 515
rect 105 505 125 525
rect 0 465 20 505
rect 105 485 150 505
rect 130 465 150 485
rect 215 465 235 590
rect 280 465 300 700
rect 320 670 360 680
rect 320 600 330 670
rect 350 600 360 670
rect 320 590 360 600
rect 385 670 425 680
rect 385 600 395 670
rect 415 600 425 670
rect 385 590 425 600
rect 340 525 360 590
rect 340 515 380 525
rect 340 495 350 515
rect 370 495 380 515
rect 340 485 380 495
rect 405 465 425 590
rect -65 455 -25 465
rect -65 385 -55 455
rect -35 385 -25 455
rect -65 375 -25 385
rect 0 455 40 465
rect 0 385 10 455
rect 30 385 40 455
rect 0 375 40 385
rect 65 455 105 465
rect 65 385 75 455
rect 95 385 105 455
rect 65 375 105 385
rect 130 455 170 465
rect 130 385 140 455
rect 160 385 170 455
rect 130 375 170 385
rect 215 455 255 465
rect 215 385 225 455
rect 245 385 255 455
rect 280 455 360 465
rect 280 445 330 455
rect 215 375 255 385
rect 320 385 330 445
rect 350 385 360 455
rect 320 375 360 385
rect 385 455 425 465
rect 385 385 395 455
rect 415 385 425 455
rect 385 375 425 385
rect -45 355 -25 375
rect 65 355 85 375
rect -45 335 85 355
rect 130 355 150 375
rect 340 355 360 375
rect 130 345 275 355
rect 130 335 245 345
rect -45 300 -5 310
rect -45 290 -35 300
rect -80 280 -35 290
rect -15 280 -5 300
rect 130 290 150 335
rect 235 325 245 335
rect 265 325 275 345
rect 340 335 425 355
rect 235 315 275 325
rect 405 290 425 335
rect -80 270 -5 280
rect 60 270 150 290
rect 210 270 340 290
rect 60 245 80 270
rect 210 245 230 270
rect 320 245 340 270
rect 405 270 455 290
rect 405 245 425 270
rect -65 235 -25 245
rect -65 165 -55 235
rect -35 165 -25 235
rect 40 235 80 245
rect 40 175 50 235
rect -65 155 -25 165
rect 0 165 50 175
rect 70 165 80 235
rect 0 155 80 165
rect 105 235 145 245
rect 105 165 115 235
rect 135 165 145 235
rect 105 155 145 165
rect 190 235 230 245
rect 190 165 200 235
rect 220 165 230 235
rect 190 155 230 165
rect 255 235 295 245
rect 255 165 265 235
rect 285 165 295 235
rect 255 155 295 165
rect 320 235 360 245
rect 320 165 330 235
rect 350 165 360 235
rect 320 155 360 165
rect 385 235 425 245
rect 385 165 395 235
rect 415 165 425 235
rect 385 155 425 165
rect -65 30 -45 155
rect -65 20 -25 30
rect -65 -50 -55 20
rect -35 -50 -25 20
rect -65 -60 -25 -50
rect 0 -80 20 155
rect 60 125 100 135
rect 60 105 70 125
rect 90 105 100 125
rect 60 95 100 105
rect 60 30 80 95
rect 125 30 145 155
rect 255 115 275 155
rect 385 135 405 155
rect 360 115 405 135
rect 190 105 280 115
rect 190 85 200 105
rect 270 85 280 105
rect 360 90 380 115
rect 190 75 280 85
rect 340 80 380 90
rect 255 30 275 75
rect 340 60 350 80
rect 370 60 380 80
rect 340 50 380 60
rect 405 75 445 85
rect 405 55 415 75
rect 435 55 445 75
rect 405 45 445 55
rect 405 30 425 45
rect 40 20 80 30
rect 40 -50 50 20
rect 70 -50 80 20
rect 40 -60 80 -50
rect 105 20 145 30
rect 105 -50 115 20
rect 135 -50 145 20
rect 105 -60 145 -50
rect 190 20 230 30
rect 190 -50 200 20
rect 220 -50 230 20
rect 190 -60 230 -50
rect 255 20 295 30
rect 255 -50 265 20
rect 285 -50 295 20
rect 255 -60 295 -50
rect 320 20 360 30
rect 320 -50 330 20
rect 350 -50 360 20
rect 320 -60 360 -50
rect 385 20 425 30
rect 385 -50 395 20
rect 415 -50 425 20
rect 385 -60 425 -50
rect 210 -80 230 -60
rect 320 -80 340 -60
rect 0 -90 100 -80
rect 0 -100 70 -90
rect 60 -110 70 -100
rect 90 -110 100 -90
rect 210 -100 340 -80
rect 60 -120 100 -110
rect -5 -130 35 -120
rect -5 -150 5 -130
rect 25 -150 35 -130
rect -5 -160 35 -150
rect 340 -130 380 -120
rect 340 -150 350 -130
rect 370 -150 380 -130
rect 340 -160 380 -150
<< viali >>
rect 10 600 30 670
rect 225 600 245 670
rect 10 385 30 455
rect 225 385 245 455
rect -55 165 -35 235
rect 200 165 220 235
rect -55 -50 -35 20
rect 200 85 270 105
rect 200 -50 220 20
rect 5 -150 25 -130
rect 350 -150 370 -130
<< metal1 >>
rect -80 670 455 685
rect -80 600 10 670
rect 30 600 225 670
rect 245 600 455 670
rect -80 455 455 600
rect -80 385 10 455
rect 30 385 225 455
rect 245 385 455 455
rect -80 370 455 385
rect -80 235 455 250
rect -80 165 -55 235
rect -35 165 200 235
rect 220 165 455 235
rect -80 105 455 165
rect -80 85 200 105
rect 270 85 455 105
rect -80 20 455 85
rect -80 -50 -55 20
rect -35 -50 200 20
rect 220 -50 455 20
rect -80 -65 455 -50
rect -80 -130 455 -120
rect -80 -150 5 -130
rect 25 -150 350 -130
rect 370 -150 455 -130
rect -80 -160 455 -150
<< end >>
